module BF( // @[:@3.2]
  input  [9:0] io_in1_re, // @[:@6.4]
  input  [9:0] io_in1_im, // @[:@6.4]
  input  [9:0] io_in2_re, // @[:@6.4]
  input  [9:0] io_in2_im, // @[:@6.4]
  output [9:0] io_out1_re, // @[:@6.4]
  output [9:0] io_out1_im, // @[:@6.4]
  output [9:0] io_out2_re, // @[:@6.4]
  output [9:0] io_out2_im // @[:@6.4]
);
  wire [10:0] _T_13; // @[R2MDC.scala 26:27:@8.4]
  wire [9:0] _T_14; // @[R2MDC.scala 26:27:@9.4]
  wire [10:0] _T_16; // @[R2MDC.scala 27:27:@12.4]
  wire [9:0] _T_17; // @[R2MDC.scala 27:27:@13.4]
  wire [10:0] _T_19; // @[R2MDC.scala 28:27:@16.4]
  wire [9:0] _T_20; // @[R2MDC.scala 28:27:@17.4]
  wire [10:0] _T_22; // @[R2MDC.scala 29:27:@20.4]
  wire [9:0] _T_23; // @[R2MDC.scala 29:27:@21.4]
  assign _T_13 = $signed(io_in1_re) + $signed(io_in2_re); // @[R2MDC.scala 26:27:@8.4]
  assign _T_14 = _T_13[9:0]; // @[R2MDC.scala 26:27:@9.4]
  assign _T_16 = $signed(io_in1_im) + $signed(io_in2_im); // @[R2MDC.scala 27:27:@12.4]
  assign _T_17 = _T_16[9:0]; // @[R2MDC.scala 27:27:@13.4]
  assign _T_19 = $signed(io_in1_re) - $signed(io_in2_re); // @[R2MDC.scala 28:27:@16.4]
  assign _T_20 = _T_19[9:0]; // @[R2MDC.scala 28:27:@17.4]
  assign _T_22 = $signed(io_in1_im) - $signed(io_in2_im); // @[R2MDC.scala 29:27:@20.4]
  assign _T_23 = _T_22[9:0]; // @[R2MDC.scala 29:27:@21.4]
  assign io_out1_re = $signed(_T_14); // @[R2MDC.scala 26:14:@11.4]
  assign io_out1_im = $signed(_T_17); // @[R2MDC.scala 27:14:@15.4]
  assign io_out2_re = $signed(_T_20); // @[R2MDC.scala 28:14:@19.4]
  assign io_out2_im = $signed(_T_23); // @[R2MDC.scala 29:14:@23.4]
endmodule
module complexMul( // @[:@25.2]
  input  [9:0] io_in1_re, // @[:@28.4]
  input  [9:0] io_in1_im, // @[:@28.4]
  input  [9:0] io_in2_re, // @[:@28.4]
  input  [9:0] io_in2_im, // @[:@28.4]
  output [9:0] io_out_re, // @[:@28.4]
  output [9:0] io_out_im // @[:@28.4]
);
  wire [10:0] _T_11; // @[R2MDC.scala 48:37:@30.4]
  wire [9:0] _T_12; // @[R2MDC.scala 48:37:@31.4]
  wire [9:0] _T_13; // @[R2MDC.scala 48:37:@32.4]
  wire [19:0] _T_14; // @[R2MDC.scala 48:24:@33.4]
  wire [10:0] _T_15; // @[R2MDC.scala 49:37:@34.4]
  wire [9:0] _T_16; // @[R2MDC.scala 49:37:@35.4]
  wire [9:0] _T_17; // @[R2MDC.scala 49:37:@36.4]
  wire [19:0] _T_18; // @[R2MDC.scala 49:24:@37.4]
  wire [10:0] _T_19; // @[R2MDC.scala 50:37:@38.4]
  wire [9:0] _T_20; // @[R2MDC.scala 50:37:@39.4]
  wire [9:0] _T_21; // @[R2MDC.scala 50:37:@40.4]
  wire [19:0] _T_22; // @[R2MDC.scala 50:24:@41.4]
  wire [20:0] _T_23; // @[R2MDC.scala 51:22:@42.4]
  wire [19:0] _T_24; // @[R2MDC.scala 51:22:@43.4]
  wire [19:0] _T_25; // @[R2MDC.scala 51:22:@44.4]
  wire [11:0] _T_26; // @[R2MDC.scala 51:28:@45.4]
  wire [20:0] _T_27; // @[R2MDC.scala 52:22:@47.4]
  wire [19:0] _T_28; // @[R2MDC.scala 52:22:@48.4]
  wire [19:0] _T_29; // @[R2MDC.scala 52:22:@49.4]
  wire [11:0] _T_30; // @[R2MDC.scala 52:28:@50.4]
  wire [9:0] _GEN_0; // @[R2MDC.scala 51:15:@46.4]
  wire [9:0] _GEN_1; // @[R2MDC.scala 52:15:@51.4]
  assign _T_11 = $signed(io_in1_re) + $signed(io_in1_im); // @[R2MDC.scala 48:37:@30.4]
  assign _T_12 = _T_11[9:0]; // @[R2MDC.scala 48:37:@31.4]
  assign _T_13 = $signed(_T_12); // @[R2MDC.scala 48:37:@32.4]
  assign _T_14 = $signed(io_in2_re) * $signed(_T_13); // @[R2MDC.scala 48:24:@33.4]
  assign _T_15 = $signed(io_in2_im) - $signed(io_in2_re); // @[R2MDC.scala 49:37:@34.4]
  assign _T_16 = _T_15[9:0]; // @[R2MDC.scala 49:37:@35.4]
  assign _T_17 = $signed(_T_16); // @[R2MDC.scala 49:37:@36.4]
  assign _T_18 = $signed(io_in1_re) * $signed(_T_17); // @[R2MDC.scala 49:24:@37.4]
  assign _T_19 = $signed(io_in2_re) + $signed(io_in2_im); // @[R2MDC.scala 50:37:@38.4]
  assign _T_20 = _T_19[9:0]; // @[R2MDC.scala 50:37:@39.4]
  assign _T_21 = $signed(_T_20); // @[R2MDC.scala 50:37:@40.4]
  assign _T_22 = $signed(io_in1_im) * $signed(_T_21); // @[R2MDC.scala 50:24:@41.4]
  assign _T_23 = $signed(_T_14) - $signed(_T_22); // @[R2MDC.scala 51:22:@42.4]
  assign _T_24 = _T_23[19:0]; // @[R2MDC.scala 51:22:@43.4]
  assign _T_25 = $signed(_T_24); // @[R2MDC.scala 51:22:@44.4]
  assign _T_26 = _T_25[19:8]; // @[R2MDC.scala 51:28:@45.4]
  assign _T_27 = $signed(_T_14) + $signed(_T_18); // @[R2MDC.scala 52:22:@47.4]
  assign _T_28 = _T_27[19:0]; // @[R2MDC.scala 52:22:@48.4]
  assign _T_29 = $signed(_T_28); // @[R2MDC.scala 52:22:@49.4]
  assign _T_30 = _T_29[19:8]; // @[R2MDC.scala 52:28:@50.4]
  assign _GEN_0 = _T_26[9:0]; // @[R2MDC.scala 51:15:@46.4]
  assign io_out_re = $signed(_GEN_0); // @[R2MDC.scala 51:15:@46.4]
  assign _GEN_1 = _T_30[9:0]; // @[R2MDC.scala 52:15:@51.4]
  assign io_out_im = $signed(_GEN_1); // @[R2MDC.scala 52:15:@51.4]
endmodule
module Switch( // @[:@53.2]
  input  [9:0] io_in1_re, // @[:@56.4]
  input  [9:0] io_in1_im, // @[:@56.4]
  input  [9:0] io_in2_re, // @[:@56.4]
  input  [9:0] io_in2_im, // @[:@56.4]
  input        io_sel, // @[:@56.4]
  output [9:0] io_out1_re, // @[:@56.4]
  output [9:0] io_out1_im, // @[:@56.4]
  output [9:0] io_out2_re, // @[:@56.4]
  output [9:0] io_out2_im // @[:@56.4]
);
  assign io_out1_re = io_sel ? $signed(io_in2_re) : $signed(io_in1_re); // @[R2MDC.scala 75:11:@60.4]
  assign io_out1_im = io_sel ? $signed(io_in2_im) : $signed(io_in1_im); // @[R2MDC.scala 75:11:@59.4]
  assign io_out2_re = io_sel ? $signed(io_in1_re) : $signed(io_in2_re); // @[R2MDC.scala 76:11:@63.4]
  assign io_out2_im = io_sel ? $signed(io_in1_im) : $signed(io_in2_im); // @[R2MDC.scala 76:11:@62.4]
endmodule
module R2MDC( // @[:@335.2]
  input        clock, // @[:@336.4]
  input        reset, // @[:@337.4]
  input  [9:0] io_dIn_re, // @[:@338.4]
  input  [9:0] io_dIn_im, // @[:@338.4]
  input        io_din_valid, // @[:@338.4]
  output [9:0] io_dOut1_re, // @[:@338.4]
  output [9:0] io_dOut1_im, // @[:@338.4]
  output [9:0] io_dOut2_re, // @[:@338.4]
  output [9:0] io_dOut2_im, // @[:@338.4]
  output       io_dout_valid // @[:@338.4]
);
  wire [9:0] BF_io_in1_re; // @[R2MDC.scala 33:22:@652.4]
  wire [9:0] BF_io_in1_im; // @[R2MDC.scala 33:22:@652.4]
  wire [9:0] BF_io_in2_re; // @[R2MDC.scala 33:22:@652.4]
  wire [9:0] BF_io_in2_im; // @[R2MDC.scala 33:22:@652.4]
  wire [9:0] BF_io_out1_re; // @[R2MDC.scala 33:22:@652.4]
  wire [9:0] BF_io_out1_im; // @[R2MDC.scala 33:22:@652.4]
  wire [9:0] BF_io_out2_re; // @[R2MDC.scala 33:22:@652.4]
  wire [9:0] BF_io_out2_im; // @[R2MDC.scala 33:22:@652.4]
  wire [9:0] complexMul_io_in1_re; // @[R2MDC.scala 60:22:@729.4]
  wire [9:0] complexMul_io_in1_im; // @[R2MDC.scala 60:22:@729.4]
  wire [9:0] complexMul_io_in2_re; // @[R2MDC.scala 60:22:@729.4]
  wire [9:0] complexMul_io_in2_im; // @[R2MDC.scala 60:22:@729.4]
  wire [9:0] complexMul_io_out_re; // @[R2MDC.scala 60:22:@729.4]
  wire [9:0] complexMul_io_out_im; // @[R2MDC.scala 60:22:@729.4]
  wire [9:0] Switch_io_in1_re; // @[R2MDC.scala 80:22:@817.4]
  wire [9:0] Switch_io_in1_im; // @[R2MDC.scala 80:22:@817.4]
  wire [9:0] Switch_io_in2_re; // @[R2MDC.scala 80:22:@817.4]
  wire [9:0] Switch_io_in2_im; // @[R2MDC.scala 80:22:@817.4]
  wire  Switch_io_sel; // @[R2MDC.scala 80:22:@817.4]
  wire [9:0] Switch_io_out1_re; // @[R2MDC.scala 80:22:@817.4]
  wire [9:0] Switch_io_out1_im; // @[R2MDC.scala 80:22:@817.4]
  wire [9:0] Switch_io_out2_re; // @[R2MDC.scala 80:22:@817.4]
  wire [9:0] Switch_io_out2_im; // @[R2MDC.scala 80:22:@817.4]
  wire [9:0] BF_1_io_in1_re; // @[R2MDC.scala 33:22:@909.4]
  wire [9:0] BF_1_io_in1_im; // @[R2MDC.scala 33:22:@909.4]
  wire [9:0] BF_1_io_in2_re; // @[R2MDC.scala 33:22:@909.4]
  wire [9:0] BF_1_io_in2_im; // @[R2MDC.scala 33:22:@909.4]
  wire [9:0] BF_1_io_out1_re; // @[R2MDC.scala 33:22:@909.4]
  wire [9:0] BF_1_io_out1_im; // @[R2MDC.scala 33:22:@909.4]
  wire [9:0] BF_1_io_out2_re; // @[R2MDC.scala 33:22:@909.4]
  wire [9:0] BF_1_io_out2_im; // @[R2MDC.scala 33:22:@909.4]
  wire [9:0] complexMul_1_io_in1_re; // @[R2MDC.scala 60:22:@954.4]
  wire [9:0] complexMul_1_io_in1_im; // @[R2MDC.scala 60:22:@954.4]
  wire [9:0] complexMul_1_io_in2_re; // @[R2MDC.scala 60:22:@954.4]
  wire [9:0] complexMul_1_io_in2_im; // @[R2MDC.scala 60:22:@954.4]
  wire [9:0] complexMul_1_io_out_re; // @[R2MDC.scala 60:22:@954.4]
  wire [9:0] complexMul_1_io_out_im; // @[R2MDC.scala 60:22:@954.4]
  wire [9:0] Switch_1_io_in1_re; // @[R2MDC.scala 80:22:@1002.4]
  wire [9:0] Switch_1_io_in1_im; // @[R2MDC.scala 80:22:@1002.4]
  wire [9:0] Switch_1_io_in2_re; // @[R2MDC.scala 80:22:@1002.4]
  wire [9:0] Switch_1_io_in2_im; // @[R2MDC.scala 80:22:@1002.4]
  wire  Switch_1_io_sel; // @[R2MDC.scala 80:22:@1002.4]
  wire [9:0] Switch_1_io_out1_re; // @[R2MDC.scala 80:22:@1002.4]
  wire [9:0] Switch_1_io_out1_im; // @[R2MDC.scala 80:22:@1002.4]
  wire [9:0] Switch_1_io_out2_re; // @[R2MDC.scala 80:22:@1002.4]
  wire [9:0] Switch_1_io_out2_im; // @[R2MDC.scala 80:22:@1002.4]
  wire [9:0] BF_2_io_in1_re; // @[R2MDC.scala 33:22:@1054.4]
  wire [9:0] BF_2_io_in1_im; // @[R2MDC.scala 33:22:@1054.4]
  wire [9:0] BF_2_io_in2_re; // @[R2MDC.scala 33:22:@1054.4]
  wire [9:0] BF_2_io_in2_im; // @[R2MDC.scala 33:22:@1054.4]
  wire [9:0] BF_2_io_out1_re; // @[R2MDC.scala 33:22:@1054.4]
  wire [9:0] BF_2_io_out1_im; // @[R2MDC.scala 33:22:@1054.4]
  wire [9:0] BF_2_io_out2_re; // @[R2MDC.scala 33:22:@1054.4]
  wire [9:0] BF_2_io_out2_im; // @[R2MDC.scala 33:22:@1054.4]
  wire [9:0] complexMul_2_io_in1_re; // @[R2MDC.scala 60:22:@1083.4]
  wire [9:0] complexMul_2_io_in1_im; // @[R2MDC.scala 60:22:@1083.4]
  wire [9:0] complexMul_2_io_in2_re; // @[R2MDC.scala 60:22:@1083.4]
  wire [9:0] complexMul_2_io_in2_im; // @[R2MDC.scala 60:22:@1083.4]
  wire [9:0] complexMul_2_io_out_re; // @[R2MDC.scala 60:22:@1083.4]
  wire [9:0] complexMul_2_io_out_im; // @[R2MDC.scala 60:22:@1083.4]
  wire [9:0] Switch_2_io_in1_re; // @[R2MDC.scala 80:22:@1111.4]
  wire [9:0] Switch_2_io_in1_im; // @[R2MDC.scala 80:22:@1111.4]
  wire [9:0] Switch_2_io_in2_re; // @[R2MDC.scala 80:22:@1111.4]
  wire [9:0] Switch_2_io_in2_im; // @[R2MDC.scala 80:22:@1111.4]
  wire  Switch_2_io_sel; // @[R2MDC.scala 80:22:@1111.4]
  wire [9:0] Switch_2_io_out1_re; // @[R2MDC.scala 80:22:@1111.4]
  wire [9:0] Switch_2_io_out1_im; // @[R2MDC.scala 80:22:@1111.4]
  wire [9:0] Switch_2_io_out2_re; // @[R2MDC.scala 80:22:@1111.4]
  wire [9:0] Switch_2_io_out2_im; // @[R2MDC.scala 80:22:@1111.4]
  wire [9:0] BF_3_io_in1_re; // @[R2MDC.scala 33:22:@1143.4]
  wire [9:0] BF_3_io_in1_im; // @[R2MDC.scala 33:22:@1143.4]
  wire [9:0] BF_3_io_in2_re; // @[R2MDC.scala 33:22:@1143.4]
  wire [9:0] BF_3_io_in2_im; // @[R2MDC.scala 33:22:@1143.4]
  wire [9:0] BF_3_io_out1_re; // @[R2MDC.scala 33:22:@1143.4]
  wire [9:0] BF_3_io_out1_im; // @[R2MDC.scala 33:22:@1143.4]
  wire [9:0] BF_3_io_out2_re; // @[R2MDC.scala 33:22:@1143.4]
  wire [9:0] BF_3_io_out2_im; // @[R2MDC.scala 33:22:@1143.4]
  wire [9:0] complexMul_3_io_in1_re; // @[R2MDC.scala 60:22:@1164.4]
  wire [9:0] complexMul_3_io_in1_im; // @[R2MDC.scala 60:22:@1164.4]
  wire [9:0] complexMul_3_io_in2_re; // @[R2MDC.scala 60:22:@1164.4]
  wire [9:0] complexMul_3_io_in2_im; // @[R2MDC.scala 60:22:@1164.4]
  wire [9:0] complexMul_3_io_out_re; // @[R2MDC.scala 60:22:@1164.4]
  wire [9:0] complexMul_3_io_out_im; // @[R2MDC.scala 60:22:@1164.4]
  wire [9:0] Switch_3_io_in1_re; // @[R2MDC.scala 80:22:@1182.4]
  wire [9:0] Switch_3_io_in1_im; // @[R2MDC.scala 80:22:@1182.4]
  wire [9:0] Switch_3_io_in2_re; // @[R2MDC.scala 80:22:@1182.4]
  wire [9:0] Switch_3_io_in2_im; // @[R2MDC.scala 80:22:@1182.4]
  wire  Switch_3_io_sel; // @[R2MDC.scala 80:22:@1182.4]
  wire [9:0] Switch_3_io_out1_re; // @[R2MDC.scala 80:22:@1182.4]
  wire [9:0] Switch_3_io_out1_im; // @[R2MDC.scala 80:22:@1182.4]
  wire [9:0] Switch_3_io_out2_re; // @[R2MDC.scala 80:22:@1182.4]
  wire [9:0] Switch_3_io_out2_im; // @[R2MDC.scala 80:22:@1182.4]
  wire [9:0] BF_4_io_in1_re; // @[R2MDC.scala 33:22:@1204.4]
  wire [9:0] BF_4_io_in1_im; // @[R2MDC.scala 33:22:@1204.4]
  wire [9:0] BF_4_io_in2_re; // @[R2MDC.scala 33:22:@1204.4]
  wire [9:0] BF_4_io_in2_im; // @[R2MDC.scala 33:22:@1204.4]
  wire [9:0] BF_4_io_out1_re; // @[R2MDC.scala 33:22:@1204.4]
  wire [9:0] BF_4_io_out1_im; // @[R2MDC.scala 33:22:@1204.4]
  wire [9:0] BF_4_io_out2_re; // @[R2MDC.scala 33:22:@1204.4]
  wire [9:0] BF_4_io_out2_im; // @[R2MDC.scala 33:22:@1204.4]
  wire [9:0] complexMul_4_io_in1_re; // @[R2MDC.scala 60:22:@1221.4]
  wire [9:0] complexMul_4_io_in1_im; // @[R2MDC.scala 60:22:@1221.4]
  wire [9:0] complexMul_4_io_in2_re; // @[R2MDC.scala 60:22:@1221.4]
  wire [9:0] complexMul_4_io_in2_im; // @[R2MDC.scala 60:22:@1221.4]
  wire [9:0] complexMul_4_io_out_re; // @[R2MDC.scala 60:22:@1221.4]
  wire [9:0] complexMul_4_io_out_im; // @[R2MDC.scala 60:22:@1221.4]
  wire [9:0] Switch_4_io_in1_re; // @[R2MDC.scala 80:22:@1234.4]
  wire [9:0] Switch_4_io_in1_im; // @[R2MDC.scala 80:22:@1234.4]
  wire [9:0] Switch_4_io_in2_re; // @[R2MDC.scala 80:22:@1234.4]
  wire [9:0] Switch_4_io_in2_im; // @[R2MDC.scala 80:22:@1234.4]
  wire  Switch_4_io_sel; // @[R2MDC.scala 80:22:@1234.4]
  wire [9:0] Switch_4_io_out1_re; // @[R2MDC.scala 80:22:@1234.4]
  wire [9:0] Switch_4_io_out1_im; // @[R2MDC.scala 80:22:@1234.4]
  wire [9:0] Switch_4_io_out2_re; // @[R2MDC.scala 80:22:@1234.4]
  wire [9:0] Switch_4_io_out2_im; // @[R2MDC.scala 80:22:@1234.4]
  wire [9:0] BF_5_io_in1_re; // @[R2MDC.scala 33:22:@1251.4]
  wire [9:0] BF_5_io_in1_im; // @[R2MDC.scala 33:22:@1251.4]
  wire [9:0] BF_5_io_in2_re; // @[R2MDC.scala 33:22:@1251.4]
  wire [9:0] BF_5_io_in2_im; // @[R2MDC.scala 33:22:@1251.4]
  wire [9:0] BF_5_io_out1_re; // @[R2MDC.scala 33:22:@1251.4]
  wire [9:0] BF_5_io_out1_im; // @[R2MDC.scala 33:22:@1251.4]
  wire [9:0] BF_5_io_out2_re; // @[R2MDC.scala 33:22:@1251.4]
  wire [9:0] BF_5_io_out2_im; // @[R2MDC.scala 33:22:@1251.4]
  reg [5:0] cnt; // @[R2MDC.scala 120:20:@340.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_18; // @[R2MDC.scala 122:16:@342.6]
  wire [5:0] _T_19; // @[R2MDC.scala 122:16:@343.6]
  wire [5:0] _GEN_0; // @[R2MDC.scala 121:21:@341.4]
  reg [9:0] _T_176_re; // @[Reg.scala 11:16:@492.4]
  reg [31:0] _RAND_1;
  reg [9:0] _T_176_im; // @[Reg.scala 11:16:@492.4]
  reg [31:0] _RAND_2;
  reg [9:0] _T_178_re; // @[Reg.scala 11:16:@497.4]
  reg [31:0] _RAND_3;
  reg [9:0] _T_178_im; // @[Reg.scala 11:16:@497.4]
  reg [31:0] _RAND_4;
  reg [9:0] _T_180_re; // @[Reg.scala 11:16:@502.4]
  reg [31:0] _RAND_5;
  reg [9:0] _T_180_im; // @[Reg.scala 11:16:@502.4]
  reg [31:0] _RAND_6;
  reg [9:0] _T_182_re; // @[Reg.scala 11:16:@507.4]
  reg [31:0] _RAND_7;
  reg [9:0] _T_182_im; // @[Reg.scala 11:16:@507.4]
  reg [31:0] _RAND_8;
  reg [9:0] _T_184_re; // @[Reg.scala 11:16:@512.4]
  reg [31:0] _RAND_9;
  reg [9:0] _T_184_im; // @[Reg.scala 11:16:@512.4]
  reg [31:0] _RAND_10;
  reg [9:0] _T_186_re; // @[Reg.scala 11:16:@517.4]
  reg [31:0] _RAND_11;
  reg [9:0] _T_186_im; // @[Reg.scala 11:16:@517.4]
  reg [31:0] _RAND_12;
  reg [9:0] _T_188_re; // @[Reg.scala 11:16:@522.4]
  reg [31:0] _RAND_13;
  reg [9:0] _T_188_im; // @[Reg.scala 11:16:@522.4]
  reg [31:0] _RAND_14;
  reg [9:0] _T_190_re; // @[Reg.scala 11:16:@527.4]
  reg [31:0] _RAND_15;
  reg [9:0] _T_190_im; // @[Reg.scala 11:16:@527.4]
  reg [31:0] _RAND_16;
  reg [9:0] _T_192_re; // @[Reg.scala 11:16:@532.4]
  reg [31:0] _RAND_17;
  reg [9:0] _T_192_im; // @[Reg.scala 11:16:@532.4]
  reg [31:0] _RAND_18;
  reg [9:0] _T_194_re; // @[Reg.scala 11:16:@537.4]
  reg [31:0] _RAND_19;
  reg [9:0] _T_194_im; // @[Reg.scala 11:16:@537.4]
  reg [31:0] _RAND_20;
  reg [9:0] _T_196_re; // @[Reg.scala 11:16:@542.4]
  reg [31:0] _RAND_21;
  reg [9:0] _T_196_im; // @[Reg.scala 11:16:@542.4]
  reg [31:0] _RAND_22;
  reg [9:0] _T_198_re; // @[Reg.scala 11:16:@547.4]
  reg [31:0] _RAND_23;
  reg [9:0] _T_198_im; // @[Reg.scala 11:16:@547.4]
  reg [31:0] _RAND_24;
  reg [9:0] _T_200_re; // @[Reg.scala 11:16:@552.4]
  reg [31:0] _RAND_25;
  reg [9:0] _T_200_im; // @[Reg.scala 11:16:@552.4]
  reg [31:0] _RAND_26;
  reg [9:0] _T_202_re; // @[Reg.scala 11:16:@557.4]
  reg [31:0] _RAND_27;
  reg [9:0] _T_202_im; // @[Reg.scala 11:16:@557.4]
  reg [31:0] _RAND_28;
  reg [9:0] _T_204_re; // @[Reg.scala 11:16:@562.4]
  reg [31:0] _RAND_29;
  reg [9:0] _T_204_im; // @[Reg.scala 11:16:@562.4]
  reg [31:0] _RAND_30;
  reg [9:0] _T_206_re; // @[Reg.scala 11:16:@567.4]
  reg [31:0] _RAND_31;
  reg [9:0] _T_206_im; // @[Reg.scala 11:16:@567.4]
  reg [31:0] _RAND_32;
  reg [9:0] _T_208_re; // @[Reg.scala 11:16:@572.4]
  reg [31:0] _RAND_33;
  reg [9:0] _T_208_im; // @[Reg.scala 11:16:@572.4]
  reg [31:0] _RAND_34;
  reg [9:0] _T_210_re; // @[Reg.scala 11:16:@577.4]
  reg [31:0] _RAND_35;
  reg [9:0] _T_210_im; // @[Reg.scala 11:16:@577.4]
  reg [31:0] _RAND_36;
  reg [9:0] _T_212_re; // @[Reg.scala 11:16:@582.4]
  reg [31:0] _RAND_37;
  reg [9:0] _T_212_im; // @[Reg.scala 11:16:@582.4]
  reg [31:0] _RAND_38;
  reg [9:0] _T_214_re; // @[Reg.scala 11:16:@587.4]
  reg [31:0] _RAND_39;
  reg [9:0] _T_214_im; // @[Reg.scala 11:16:@587.4]
  reg [31:0] _RAND_40;
  reg [9:0] _T_216_re; // @[Reg.scala 11:16:@592.4]
  reg [31:0] _RAND_41;
  reg [9:0] _T_216_im; // @[Reg.scala 11:16:@592.4]
  reg [31:0] _RAND_42;
  reg [9:0] _T_218_re; // @[Reg.scala 11:16:@597.4]
  reg [31:0] _RAND_43;
  reg [9:0] _T_218_im; // @[Reg.scala 11:16:@597.4]
  reg [31:0] _RAND_44;
  reg [9:0] _T_220_re; // @[Reg.scala 11:16:@602.4]
  reg [31:0] _RAND_45;
  reg [9:0] _T_220_im; // @[Reg.scala 11:16:@602.4]
  reg [31:0] _RAND_46;
  reg [9:0] _T_222_re; // @[Reg.scala 11:16:@607.4]
  reg [31:0] _RAND_47;
  reg [9:0] _T_222_im; // @[Reg.scala 11:16:@607.4]
  reg [31:0] _RAND_48;
  reg [9:0] _T_224_re; // @[Reg.scala 11:16:@612.4]
  reg [31:0] _RAND_49;
  reg [9:0] _T_224_im; // @[Reg.scala 11:16:@612.4]
  reg [31:0] _RAND_50;
  reg [9:0] _T_226_re; // @[Reg.scala 11:16:@617.4]
  reg [31:0] _RAND_51;
  reg [9:0] _T_226_im; // @[Reg.scala 11:16:@617.4]
  reg [31:0] _RAND_52;
  reg [9:0] _T_228_re; // @[Reg.scala 11:16:@622.4]
  reg [31:0] _RAND_53;
  reg [9:0] _T_228_im; // @[Reg.scala 11:16:@622.4]
  reg [31:0] _RAND_54;
  reg [9:0] _T_230_re; // @[Reg.scala 11:16:@627.4]
  reg [31:0] _RAND_55;
  reg [9:0] _T_230_im; // @[Reg.scala 11:16:@627.4]
  reg [31:0] _RAND_56;
  reg [9:0] _T_232_re; // @[Reg.scala 11:16:@632.4]
  reg [31:0] _RAND_57;
  reg [9:0] _T_232_im; // @[Reg.scala 11:16:@632.4]
  reg [31:0] _RAND_58;
  reg [9:0] _T_234_re; // @[Reg.scala 11:16:@637.4]
  reg [31:0] _RAND_59;
  reg [9:0] _T_234_im; // @[Reg.scala 11:16:@637.4]
  reg [31:0] _RAND_60;
  reg [9:0] _T_236_re; // @[Reg.scala 11:16:@642.4]
  reg [31:0] _RAND_61;
  reg [9:0] _T_236_im; // @[Reg.scala 11:16:@642.4]
  reg [31:0] _RAND_62;
  reg [9:0] _T_238_re; // @[Reg.scala 11:16:@647.4]
  reg [31:0] _RAND_63;
  reg [9:0] _T_238_im; // @[Reg.scala 11:16:@647.4]
  reg [31:0] _RAND_64;
  wire [4:0] _T_239; // @[R2MDC.scala 131:23:@659.4]
  wire [9:0] _GEN_66; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_67; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_68; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_69; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_70; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_71; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_72; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_73; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_74; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_75; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_76; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_77; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_78; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_79; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_80; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_81; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_82; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_83; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_84; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_85; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_86; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_87; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_88; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_89; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_90; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_91; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_92; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_93; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_94; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_95; // @[R2MDC.scala 115:12:@694.4]
  wire [9:0] _GEN_98; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_99; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_100; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_101; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_102; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_103; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_104; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_105; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_106; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_107; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_108; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_109; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_110; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_111; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_112; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_113; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_114; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_115; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_116; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_117; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_118; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_119; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_120; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_121; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_122; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_123; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_124; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_125; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_126; // @[R2MDC.scala 116:12:@728.4]
  wire [9:0] _GEN_127; // @[R2MDC.scala 116:12:@728.4]
  reg [9:0] _T_386_re; // @[Reg.scala 11:16:@736.4]
  reg [31:0] _RAND_65;
  reg [9:0] _T_386_im; // @[Reg.scala 11:16:@736.4]
  reg [31:0] _RAND_66;
  reg [9:0] _T_388_re; // @[Reg.scala 11:16:@741.4]
  reg [31:0] _RAND_67;
  reg [9:0] _T_388_im; // @[Reg.scala 11:16:@741.4]
  reg [31:0] _RAND_68;
  reg [9:0] _T_390_re; // @[Reg.scala 11:16:@746.4]
  reg [31:0] _RAND_69;
  reg [9:0] _T_390_im; // @[Reg.scala 11:16:@746.4]
  reg [31:0] _RAND_70;
  reg [9:0] _T_392_re; // @[Reg.scala 11:16:@751.4]
  reg [31:0] _RAND_71;
  reg [9:0] _T_392_im; // @[Reg.scala 11:16:@751.4]
  reg [31:0] _RAND_72;
  reg [9:0] _T_394_re; // @[Reg.scala 11:16:@756.4]
  reg [31:0] _RAND_73;
  reg [9:0] _T_394_im; // @[Reg.scala 11:16:@756.4]
  reg [31:0] _RAND_74;
  reg [9:0] _T_396_re; // @[Reg.scala 11:16:@761.4]
  reg [31:0] _RAND_75;
  reg [9:0] _T_396_im; // @[Reg.scala 11:16:@761.4]
  reg [31:0] _RAND_76;
  reg [9:0] _T_398_re; // @[Reg.scala 11:16:@766.4]
  reg [31:0] _RAND_77;
  reg [9:0] _T_398_im; // @[Reg.scala 11:16:@766.4]
  reg [31:0] _RAND_78;
  reg [9:0] _T_400_re; // @[Reg.scala 11:16:@771.4]
  reg [31:0] _RAND_79;
  reg [9:0] _T_400_im; // @[Reg.scala 11:16:@771.4]
  reg [31:0] _RAND_80;
  reg [9:0] _T_402_re; // @[Reg.scala 11:16:@776.4]
  reg [31:0] _RAND_81;
  reg [9:0] _T_402_im; // @[Reg.scala 11:16:@776.4]
  reg [31:0] _RAND_82;
  reg [9:0] _T_404_re; // @[Reg.scala 11:16:@781.4]
  reg [31:0] _RAND_83;
  reg [9:0] _T_404_im; // @[Reg.scala 11:16:@781.4]
  reg [31:0] _RAND_84;
  reg [9:0] _T_406_re; // @[Reg.scala 11:16:@786.4]
  reg [31:0] _RAND_85;
  reg [9:0] _T_406_im; // @[Reg.scala 11:16:@786.4]
  reg [31:0] _RAND_86;
  reg [9:0] _T_408_re; // @[Reg.scala 11:16:@791.4]
  reg [31:0] _RAND_87;
  reg [9:0] _T_408_im; // @[Reg.scala 11:16:@791.4]
  reg [31:0] _RAND_88;
  reg [9:0] _T_410_re; // @[Reg.scala 11:16:@796.4]
  reg [31:0] _RAND_89;
  reg [9:0] _T_410_im; // @[Reg.scala 11:16:@796.4]
  reg [31:0] _RAND_90;
  reg [9:0] _T_412_re; // @[Reg.scala 11:16:@801.4]
  reg [31:0] _RAND_91;
  reg [9:0] _T_412_im; // @[Reg.scala 11:16:@801.4]
  reg [31:0] _RAND_92;
  reg [9:0] _T_414_re; // @[Reg.scala 11:16:@806.4]
  reg [31:0] _RAND_93;
  reg [9:0] _T_414_im; // @[Reg.scala 11:16:@806.4]
  reg [31:0] _RAND_94;
  reg [9:0] _T_416_re; // @[Reg.scala 11:16:@811.4]
  reg [31:0] _RAND_95;
  reg [9:0] _T_416_im; // @[Reg.scala 11:16:@811.4]
  reg [31:0] _RAND_96;
  reg [9:0] _T_420_re; // @[Reg.scala 11:16:@829.4]
  reg [31:0] _RAND_97;
  reg [9:0] _T_420_im; // @[Reg.scala 11:16:@829.4]
  reg [31:0] _RAND_98;
  reg [9:0] _T_422_re; // @[Reg.scala 11:16:@834.4]
  reg [31:0] _RAND_99;
  reg [9:0] _T_422_im; // @[Reg.scala 11:16:@834.4]
  reg [31:0] _RAND_100;
  reg [9:0] _T_424_re; // @[Reg.scala 11:16:@839.4]
  reg [31:0] _RAND_101;
  reg [9:0] _T_424_im; // @[Reg.scala 11:16:@839.4]
  reg [31:0] _RAND_102;
  reg [9:0] _T_426_re; // @[Reg.scala 11:16:@844.4]
  reg [31:0] _RAND_103;
  reg [9:0] _T_426_im; // @[Reg.scala 11:16:@844.4]
  reg [31:0] _RAND_104;
  reg [9:0] _T_428_re; // @[Reg.scala 11:16:@849.4]
  reg [31:0] _RAND_105;
  reg [9:0] _T_428_im; // @[Reg.scala 11:16:@849.4]
  reg [31:0] _RAND_106;
  reg [9:0] _T_430_re; // @[Reg.scala 11:16:@854.4]
  reg [31:0] _RAND_107;
  reg [9:0] _T_430_im; // @[Reg.scala 11:16:@854.4]
  reg [31:0] _RAND_108;
  reg [9:0] _T_432_re; // @[Reg.scala 11:16:@859.4]
  reg [31:0] _RAND_109;
  reg [9:0] _T_432_im; // @[Reg.scala 11:16:@859.4]
  reg [31:0] _RAND_110;
  reg [9:0] _T_434_re; // @[Reg.scala 11:16:@864.4]
  reg [31:0] _RAND_111;
  reg [9:0] _T_434_im; // @[Reg.scala 11:16:@864.4]
  reg [31:0] _RAND_112;
  reg [9:0] _T_436_re; // @[Reg.scala 11:16:@869.4]
  reg [31:0] _RAND_113;
  reg [9:0] _T_436_im; // @[Reg.scala 11:16:@869.4]
  reg [31:0] _RAND_114;
  reg [9:0] _T_438_re; // @[Reg.scala 11:16:@874.4]
  reg [31:0] _RAND_115;
  reg [9:0] _T_438_im; // @[Reg.scala 11:16:@874.4]
  reg [31:0] _RAND_116;
  reg [9:0] _T_440_re; // @[Reg.scala 11:16:@879.4]
  reg [31:0] _RAND_117;
  reg [9:0] _T_440_im; // @[Reg.scala 11:16:@879.4]
  reg [31:0] _RAND_118;
  reg [9:0] _T_442_re; // @[Reg.scala 11:16:@884.4]
  reg [31:0] _RAND_119;
  reg [9:0] _T_442_im; // @[Reg.scala 11:16:@884.4]
  reg [31:0] _RAND_120;
  reg [9:0] _T_444_re; // @[Reg.scala 11:16:@889.4]
  reg [31:0] _RAND_121;
  reg [9:0] _T_444_im; // @[Reg.scala 11:16:@889.4]
  reg [31:0] _RAND_122;
  reg [9:0] _T_446_re; // @[Reg.scala 11:16:@894.4]
  reg [31:0] _RAND_123;
  reg [9:0] _T_446_im; // @[Reg.scala 11:16:@894.4]
  reg [31:0] _RAND_124;
  reg [9:0] _T_448_re; // @[Reg.scala 11:16:@899.4]
  reg [31:0] _RAND_125;
  reg [9:0] _T_448_im; // @[Reg.scala 11:16:@899.4]
  reg [31:0] _RAND_126;
  reg [9:0] _T_450_re; // @[Reg.scala 11:16:@904.4]
  reg [31:0] _RAND_127;
  reg [9:0] _T_450_im; // @[Reg.scala 11:16:@904.4]
  reg [31:0] _RAND_128;
  wire [3:0] _T_451; // @[R2MDC.scala 144:23:@916.4]
  wire [9:0] _GEN_194; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_195; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_196; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_197; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_198; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_199; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_200; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_201; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_202; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_203; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_204; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_205; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_206; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_207; // @[R2MDC.scala 115:12:@935.4]
  wire [9:0] _GEN_210; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_211; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_212; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_213; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_214; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_215; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_216; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_217; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_218; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_219; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_220; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_221; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_222; // @[R2MDC.scala 116:12:@953.4]
  wire [9:0] _GEN_223; // @[R2MDC.scala 116:12:@953.4]
  reg [9:0] _T_534_re; // @[Reg.scala 11:16:@961.4]
  reg [31:0] _RAND_129;
  reg [9:0] _T_534_im; // @[Reg.scala 11:16:@961.4]
  reg [31:0] _RAND_130;
  reg [9:0] _T_536_re; // @[Reg.scala 11:16:@966.4]
  reg [31:0] _RAND_131;
  reg [9:0] _T_536_im; // @[Reg.scala 11:16:@966.4]
  reg [31:0] _RAND_132;
  reg [9:0] _T_538_re; // @[Reg.scala 11:16:@971.4]
  reg [31:0] _RAND_133;
  reg [9:0] _T_538_im; // @[Reg.scala 11:16:@971.4]
  reg [31:0] _RAND_134;
  reg [9:0] _T_540_re; // @[Reg.scala 11:16:@976.4]
  reg [31:0] _RAND_135;
  reg [9:0] _T_540_im; // @[Reg.scala 11:16:@976.4]
  reg [31:0] _RAND_136;
  reg [9:0] _T_542_re; // @[Reg.scala 11:16:@981.4]
  reg [31:0] _RAND_137;
  reg [9:0] _T_542_im; // @[Reg.scala 11:16:@981.4]
  reg [31:0] _RAND_138;
  reg [9:0] _T_544_re; // @[Reg.scala 11:16:@986.4]
  reg [31:0] _RAND_139;
  reg [9:0] _T_544_im; // @[Reg.scala 11:16:@986.4]
  reg [31:0] _RAND_140;
  reg [9:0] _T_546_re; // @[Reg.scala 11:16:@991.4]
  reg [31:0] _RAND_141;
  reg [9:0] _T_546_im; // @[Reg.scala 11:16:@991.4]
  reg [31:0] _RAND_142;
  reg [9:0] _T_548_re; // @[Reg.scala 11:16:@996.4]
  reg [31:0] _RAND_143;
  reg [9:0] _T_548_im; // @[Reg.scala 11:16:@996.4]
  reg [31:0] _RAND_144;
  reg [9:0] _T_552_re; // @[Reg.scala 11:16:@1014.4]
  reg [31:0] _RAND_145;
  reg [9:0] _T_552_im; // @[Reg.scala 11:16:@1014.4]
  reg [31:0] _RAND_146;
  reg [9:0] _T_554_re; // @[Reg.scala 11:16:@1019.4]
  reg [31:0] _RAND_147;
  reg [9:0] _T_554_im; // @[Reg.scala 11:16:@1019.4]
  reg [31:0] _RAND_148;
  reg [9:0] _T_556_re; // @[Reg.scala 11:16:@1024.4]
  reg [31:0] _RAND_149;
  reg [9:0] _T_556_im; // @[Reg.scala 11:16:@1024.4]
  reg [31:0] _RAND_150;
  reg [9:0] _T_558_re; // @[Reg.scala 11:16:@1029.4]
  reg [31:0] _RAND_151;
  reg [9:0] _T_558_im; // @[Reg.scala 11:16:@1029.4]
  reg [31:0] _RAND_152;
  reg [9:0] _T_560_re; // @[Reg.scala 11:16:@1034.4]
  reg [31:0] _RAND_153;
  reg [9:0] _T_560_im; // @[Reg.scala 11:16:@1034.4]
  reg [31:0] _RAND_154;
  reg [9:0] _T_562_re; // @[Reg.scala 11:16:@1039.4]
  reg [31:0] _RAND_155;
  reg [9:0] _T_562_im; // @[Reg.scala 11:16:@1039.4]
  reg [31:0] _RAND_156;
  reg [9:0] _T_564_re; // @[Reg.scala 11:16:@1044.4]
  reg [31:0] _RAND_157;
  reg [9:0] _T_564_im; // @[Reg.scala 11:16:@1044.4]
  reg [31:0] _RAND_158;
  reg [9:0] _T_566_re; // @[Reg.scala 11:16:@1049.4]
  reg [31:0] _RAND_159;
  reg [9:0] _T_566_im; // @[Reg.scala 11:16:@1049.4]
  reg [31:0] _RAND_160;
  wire [2:0] _T_567; // @[R2MDC.scala 144:23:@1061.4]
  wire [9:0] _GEN_258; // @[R2MDC.scala 115:12:@1072.4]
  wire [9:0] _GEN_259; // @[R2MDC.scala 115:12:@1072.4]
  wire [9:0] _GEN_260; // @[R2MDC.scala 115:12:@1072.4]
  wire [9:0] _GEN_261; // @[R2MDC.scala 115:12:@1072.4]
  wire [9:0] _GEN_262; // @[R2MDC.scala 115:12:@1072.4]
  wire [9:0] _GEN_263; // @[R2MDC.scala 115:12:@1072.4]
  wire [9:0] _GEN_266; // @[R2MDC.scala 116:12:@1082.4]
  wire [9:0] _GEN_267; // @[R2MDC.scala 116:12:@1082.4]
  wire [9:0] _GEN_268; // @[R2MDC.scala 116:12:@1082.4]
  wire [9:0] _GEN_269; // @[R2MDC.scala 116:12:@1082.4]
  wire [9:0] _GEN_270; // @[R2MDC.scala 116:12:@1082.4]
  wire [9:0] _GEN_271; // @[R2MDC.scala 116:12:@1082.4]
  reg [9:0] _T_618_re; // @[Reg.scala 11:16:@1090.4]
  reg [31:0] _RAND_161;
  reg [9:0] _T_618_im; // @[Reg.scala 11:16:@1090.4]
  reg [31:0] _RAND_162;
  reg [9:0] _T_620_re; // @[Reg.scala 11:16:@1095.4]
  reg [31:0] _RAND_163;
  reg [9:0] _T_620_im; // @[Reg.scala 11:16:@1095.4]
  reg [31:0] _RAND_164;
  reg [9:0] _T_622_re; // @[Reg.scala 11:16:@1100.4]
  reg [31:0] _RAND_165;
  reg [9:0] _T_622_im; // @[Reg.scala 11:16:@1100.4]
  reg [31:0] _RAND_166;
  reg [9:0] _T_624_re; // @[Reg.scala 11:16:@1105.4]
  reg [31:0] _RAND_167;
  reg [9:0] _T_624_im; // @[Reg.scala 11:16:@1105.4]
  reg [31:0] _RAND_168;
  reg [9:0] _T_628_re; // @[Reg.scala 11:16:@1123.4]
  reg [31:0] _RAND_169;
  reg [9:0] _T_628_im; // @[Reg.scala 11:16:@1123.4]
  reg [31:0] _RAND_170;
  reg [9:0] _T_630_re; // @[Reg.scala 11:16:@1128.4]
  reg [31:0] _RAND_171;
  reg [9:0] _T_630_im; // @[Reg.scala 11:16:@1128.4]
  reg [31:0] _RAND_172;
  reg [9:0] _T_632_re; // @[Reg.scala 11:16:@1133.4]
  reg [31:0] _RAND_173;
  reg [9:0] _T_632_im; // @[Reg.scala 11:16:@1133.4]
  reg [31:0] _RAND_174;
  reg [9:0] _T_634_re; // @[Reg.scala 11:16:@1138.4]
  reg [31:0] _RAND_175;
  reg [9:0] _T_634_im; // @[Reg.scala 11:16:@1138.4]
  reg [31:0] _RAND_176;
  wire [1:0] _T_635; // @[R2MDC.scala 144:23:@1150.4]
  wire [9:0] _GEN_290; // @[R2MDC.scala 115:12:@1157.4]
  wire [9:0] _GEN_291; // @[R2MDC.scala 115:12:@1157.4]
  wire [9:0] _GEN_294; // @[R2MDC.scala 116:12:@1163.4]
  wire [9:0] _GEN_295; // @[R2MDC.scala 116:12:@1163.4]
  reg [9:0] _T_670_re; // @[Reg.scala 11:16:@1171.4]
  reg [31:0] _RAND_177;
  reg [9:0] _T_670_im; // @[Reg.scala 11:16:@1171.4]
  reg [31:0] _RAND_178;
  reg [9:0] _T_672_re; // @[Reg.scala 11:16:@1176.4]
  reg [31:0] _RAND_179;
  reg [9:0] _T_672_im; // @[Reg.scala 11:16:@1176.4]
  reg [31:0] _RAND_180;
  reg [9:0] _T_676_re; // @[Reg.scala 11:16:@1194.4]
  reg [31:0] _RAND_181;
  reg [9:0] _T_676_im; // @[Reg.scala 11:16:@1194.4]
  reg [31:0] _RAND_182;
  reg [9:0] _T_678_re; // @[Reg.scala 11:16:@1199.4]
  reg [31:0] _RAND_183;
  reg [9:0] _T_678_im; // @[Reg.scala 11:16:@1199.4]
  reg [31:0] _RAND_184;
  wire  _T_679; // @[R2MDC.scala 144:23:@1211.4]
  reg [9:0] _T_706_re; // @[Reg.scala 11:16:@1228.4]
  reg [31:0] _RAND_185;
  reg [9:0] _T_706_im; // @[Reg.scala 11:16:@1228.4]
  reg [31:0] _RAND_186;
  reg [9:0] _T_710_re; // @[Reg.scala 11:16:@1246.4]
  reg [31:0] _RAND_187;
  reg [9:0] _T_710_im; // @[Reg.scala 11:16:@1246.4]
  reg [31:0] _RAND_188;
  reg [9:0] _T_712_re; // @[R2MDC.scala 161:22:@1262.4]
  reg [31:0] _RAND_189;
  reg [9:0] _T_712_im; // @[R2MDC.scala 161:22:@1262.4]
  reg [31:0] _RAND_190;
  reg [9:0] _T_714_re; // @[R2MDC.scala 162:22:@1267.4]
  reg [31:0] _RAND_191;
  reg [9:0] _T_714_im; // @[R2MDC.scala 162:22:@1267.4]
  reg [31:0] _RAND_192;
  reg  _T_717; // @[Reg.scala 11:16:@1272.4]
  reg [31:0] _RAND_193;
  reg  _T_719; // @[Reg.scala 11:16:@1276.4]
  reg [31:0] _RAND_194;
  reg  _T_721; // @[Reg.scala 11:16:@1280.4]
  reg [31:0] _RAND_195;
  reg  _T_723; // @[Reg.scala 11:16:@1284.4]
  reg [31:0] _RAND_196;
  reg  _T_725; // @[Reg.scala 11:16:@1288.4]
  reg [31:0] _RAND_197;
  reg  _T_727; // @[Reg.scala 11:16:@1292.4]
  reg [31:0] _RAND_198;
  reg  _T_729; // @[Reg.scala 11:16:@1296.4]
  reg [31:0] _RAND_199;
  reg  _T_731; // @[Reg.scala 11:16:@1300.4]
  reg [31:0] _RAND_200;
  reg  _T_733; // @[Reg.scala 11:16:@1304.4]
  reg [31:0] _RAND_201;
  reg  _T_735; // @[Reg.scala 11:16:@1308.4]
  reg [31:0] _RAND_202;
  reg  _T_737; // @[Reg.scala 11:16:@1312.4]
  reg [31:0] _RAND_203;
  reg  _T_739; // @[Reg.scala 11:16:@1316.4]
  reg [31:0] _RAND_204;
  reg  _T_741; // @[Reg.scala 11:16:@1320.4]
  reg [31:0] _RAND_205;
  reg  _T_743; // @[Reg.scala 11:16:@1324.4]
  reg [31:0] _RAND_206;
  reg  _T_745; // @[Reg.scala 11:16:@1328.4]
  reg [31:0] _RAND_207;
  reg  _T_747; // @[Reg.scala 11:16:@1332.4]
  reg [31:0] _RAND_208;
  reg  _T_749; // @[Reg.scala 11:16:@1336.4]
  reg [31:0] _RAND_209;
  reg  _T_751; // @[Reg.scala 11:16:@1340.4]
  reg [31:0] _RAND_210;
  reg  _T_753; // @[Reg.scala 11:16:@1344.4]
  reg [31:0] _RAND_211;
  reg  _T_755; // @[Reg.scala 11:16:@1348.4]
  reg [31:0] _RAND_212;
  reg  _T_757; // @[Reg.scala 11:16:@1352.4]
  reg [31:0] _RAND_213;
  reg  _T_759; // @[Reg.scala 11:16:@1356.4]
  reg [31:0] _RAND_214;
  reg  _T_761; // @[Reg.scala 11:16:@1360.4]
  reg [31:0] _RAND_215;
  reg  _T_763; // @[Reg.scala 11:16:@1364.4]
  reg [31:0] _RAND_216;
  reg  _T_765; // @[Reg.scala 11:16:@1368.4]
  reg [31:0] _RAND_217;
  reg  _T_767; // @[Reg.scala 11:16:@1372.4]
  reg [31:0] _RAND_218;
  reg  _T_769; // @[Reg.scala 11:16:@1376.4]
  reg [31:0] _RAND_219;
  reg  _T_771; // @[Reg.scala 11:16:@1380.4]
  reg [31:0] _RAND_220;
  reg  _T_773; // @[Reg.scala 11:16:@1384.4]
  reg [31:0] _RAND_221;
  reg  _T_775; // @[Reg.scala 11:16:@1388.4]
  reg [31:0] _RAND_222;
  reg  _T_777; // @[Reg.scala 11:16:@1392.4]
  reg [31:0] _RAND_223;
  reg  _T_779; // @[Reg.scala 11:16:@1396.4]
  reg [31:0] _RAND_224;
  reg  _T_781; // @[Reg.scala 11:16:@1400.4]
  reg [31:0] _RAND_225;
  reg  _T_783; // @[Reg.scala 11:16:@1404.4]
  reg [31:0] _RAND_226;
  reg  _T_785; // @[Reg.scala 11:16:@1408.4]
  reg [31:0] _RAND_227;
  reg  _T_787; // @[Reg.scala 11:16:@1412.4]
  reg [31:0] _RAND_228;
  reg  _T_789; // @[Reg.scala 11:16:@1416.4]
  reg [31:0] _RAND_229;
  reg  _T_791; // @[Reg.scala 11:16:@1420.4]
  reg [31:0] _RAND_230;
  reg  _T_793; // @[Reg.scala 11:16:@1424.4]
  reg [31:0] _RAND_231;
  reg  _T_795; // @[Reg.scala 11:16:@1428.4]
  reg [31:0] _RAND_232;
  reg  _T_797; // @[Reg.scala 11:16:@1432.4]
  reg [31:0] _RAND_233;
  reg  _T_799; // @[Reg.scala 11:16:@1436.4]
  reg [31:0] _RAND_234;
  reg  _T_801; // @[Reg.scala 11:16:@1440.4]
  reg [31:0] _RAND_235;
  reg  _T_803; // @[Reg.scala 11:16:@1444.4]
  reg [31:0] _RAND_236;
  reg  _T_805; // @[Reg.scala 11:16:@1448.4]
  reg [31:0] _RAND_237;
  reg  _T_807; // @[Reg.scala 11:16:@1452.4]
  reg [31:0] _RAND_238;
  reg  _T_809; // @[Reg.scala 11:16:@1456.4]
  reg [31:0] _RAND_239;
  reg  _T_811; // @[Reg.scala 11:16:@1460.4]
  reg [31:0] _RAND_240;
  reg  _T_813; // @[Reg.scala 11:16:@1464.4]
  reg [31:0] _RAND_241;
  reg  _T_815; // @[Reg.scala 11:16:@1468.4]
  reg [31:0] _RAND_242;
  reg  _T_817; // @[Reg.scala 11:16:@1472.4]
  reg [31:0] _RAND_243;
  reg  _T_819; // @[Reg.scala 11:16:@1476.4]
  reg [31:0] _RAND_244;
  reg  _T_821; // @[Reg.scala 11:16:@1480.4]
  reg [31:0] _RAND_245;
  reg  _T_823; // @[Reg.scala 11:16:@1484.4]
  reg [31:0] _RAND_246;
  reg  _T_825; // @[Reg.scala 11:16:@1488.4]
  reg [31:0] _RAND_247;
  reg  _T_827; // @[Reg.scala 11:16:@1492.4]
  reg [31:0] _RAND_248;
  reg  _T_829; // @[Reg.scala 11:16:@1496.4]
  reg [31:0] _RAND_249;
  reg  _T_831; // @[Reg.scala 11:16:@1500.4]
  reg [31:0] _RAND_250;
  reg  _T_833; // @[Reg.scala 11:16:@1504.4]
  reg [31:0] _RAND_251;
  reg  _T_835; // @[Reg.scala 11:16:@1508.4]
  reg [31:0] _RAND_252;
  reg  _T_837; // @[Reg.scala 11:16:@1512.4]
  reg [31:0] _RAND_253;
  reg  _T_839; // @[Reg.scala 11:16:@1516.4]
  reg [31:0] _RAND_254;
  reg  _T_841; // @[Reg.scala 11:16:@1520.4]
  reg [31:0] _RAND_255;
  reg  _T_843; // @[Reg.scala 11:16:@1524.4]
  reg [31:0] _RAND_256;
  BF BF ( // @[R2MDC.scala 33:22:@652.4]
    .io_in1_re(BF_io_in1_re),
    .io_in1_im(BF_io_in1_im),
    .io_in2_re(BF_io_in2_re),
    .io_in2_im(BF_io_in2_im),
    .io_out1_re(BF_io_out1_re),
    .io_out1_im(BF_io_out1_im),
    .io_out2_re(BF_io_out2_re),
    .io_out2_im(BF_io_out2_im)
  );
  complexMul complexMul ( // @[R2MDC.scala 60:22:@729.4]
    .io_in1_re(complexMul_io_in1_re),
    .io_in1_im(complexMul_io_in1_im),
    .io_in2_re(complexMul_io_in2_re),
    .io_in2_im(complexMul_io_in2_im),
    .io_out_re(complexMul_io_out_re),
    .io_out_im(complexMul_io_out_im)
  );
  Switch Switch ( // @[R2MDC.scala 80:22:@817.4]
    .io_in1_re(Switch_io_in1_re),
    .io_in1_im(Switch_io_in1_im),
    .io_in2_re(Switch_io_in2_re),
    .io_in2_im(Switch_io_in2_im),
    .io_sel(Switch_io_sel),
    .io_out1_re(Switch_io_out1_re),
    .io_out1_im(Switch_io_out1_im),
    .io_out2_re(Switch_io_out2_re),
    .io_out2_im(Switch_io_out2_im)
  );
  BF BF_1 ( // @[R2MDC.scala 33:22:@909.4]
    .io_in1_re(BF_1_io_in1_re),
    .io_in1_im(BF_1_io_in1_im),
    .io_in2_re(BF_1_io_in2_re),
    .io_in2_im(BF_1_io_in2_im),
    .io_out1_re(BF_1_io_out1_re),
    .io_out1_im(BF_1_io_out1_im),
    .io_out2_re(BF_1_io_out2_re),
    .io_out2_im(BF_1_io_out2_im)
  );
  complexMul complexMul_1 ( // @[R2MDC.scala 60:22:@954.4]
    .io_in1_re(complexMul_1_io_in1_re),
    .io_in1_im(complexMul_1_io_in1_im),
    .io_in2_re(complexMul_1_io_in2_re),
    .io_in2_im(complexMul_1_io_in2_im),
    .io_out_re(complexMul_1_io_out_re),
    .io_out_im(complexMul_1_io_out_im)
  );
  Switch Switch_1 ( // @[R2MDC.scala 80:22:@1002.4]
    .io_in1_re(Switch_1_io_in1_re),
    .io_in1_im(Switch_1_io_in1_im),
    .io_in2_re(Switch_1_io_in2_re),
    .io_in2_im(Switch_1_io_in2_im),
    .io_sel(Switch_1_io_sel),
    .io_out1_re(Switch_1_io_out1_re),
    .io_out1_im(Switch_1_io_out1_im),
    .io_out2_re(Switch_1_io_out2_re),
    .io_out2_im(Switch_1_io_out2_im)
  );
  BF BF_2 ( // @[R2MDC.scala 33:22:@1054.4]
    .io_in1_re(BF_2_io_in1_re),
    .io_in1_im(BF_2_io_in1_im),
    .io_in2_re(BF_2_io_in2_re),
    .io_in2_im(BF_2_io_in2_im),
    .io_out1_re(BF_2_io_out1_re),
    .io_out1_im(BF_2_io_out1_im),
    .io_out2_re(BF_2_io_out2_re),
    .io_out2_im(BF_2_io_out2_im)
  );
  complexMul complexMul_2 ( // @[R2MDC.scala 60:22:@1083.4]
    .io_in1_re(complexMul_2_io_in1_re),
    .io_in1_im(complexMul_2_io_in1_im),
    .io_in2_re(complexMul_2_io_in2_re),
    .io_in2_im(complexMul_2_io_in2_im),
    .io_out_re(complexMul_2_io_out_re),
    .io_out_im(complexMul_2_io_out_im)
  );
  Switch Switch_2 ( // @[R2MDC.scala 80:22:@1111.4]
    .io_in1_re(Switch_2_io_in1_re),
    .io_in1_im(Switch_2_io_in1_im),
    .io_in2_re(Switch_2_io_in2_re),
    .io_in2_im(Switch_2_io_in2_im),
    .io_sel(Switch_2_io_sel),
    .io_out1_re(Switch_2_io_out1_re),
    .io_out1_im(Switch_2_io_out1_im),
    .io_out2_re(Switch_2_io_out2_re),
    .io_out2_im(Switch_2_io_out2_im)
  );
  BF BF_3 ( // @[R2MDC.scala 33:22:@1143.4]
    .io_in1_re(BF_3_io_in1_re),
    .io_in1_im(BF_3_io_in1_im),
    .io_in2_re(BF_3_io_in2_re),
    .io_in2_im(BF_3_io_in2_im),
    .io_out1_re(BF_3_io_out1_re),
    .io_out1_im(BF_3_io_out1_im),
    .io_out2_re(BF_3_io_out2_re),
    .io_out2_im(BF_3_io_out2_im)
  );
  complexMul complexMul_3 ( // @[R2MDC.scala 60:22:@1164.4]
    .io_in1_re(complexMul_3_io_in1_re),
    .io_in1_im(complexMul_3_io_in1_im),
    .io_in2_re(complexMul_3_io_in2_re),
    .io_in2_im(complexMul_3_io_in2_im),
    .io_out_re(complexMul_3_io_out_re),
    .io_out_im(complexMul_3_io_out_im)
  );
  Switch Switch_3 ( // @[R2MDC.scala 80:22:@1182.4]
    .io_in1_re(Switch_3_io_in1_re),
    .io_in1_im(Switch_3_io_in1_im),
    .io_in2_re(Switch_3_io_in2_re),
    .io_in2_im(Switch_3_io_in2_im),
    .io_sel(Switch_3_io_sel),
    .io_out1_re(Switch_3_io_out1_re),
    .io_out1_im(Switch_3_io_out1_im),
    .io_out2_re(Switch_3_io_out2_re),
    .io_out2_im(Switch_3_io_out2_im)
  );
  BF BF_4 ( // @[R2MDC.scala 33:22:@1204.4]
    .io_in1_re(BF_4_io_in1_re),
    .io_in1_im(BF_4_io_in1_im),
    .io_in2_re(BF_4_io_in2_re),
    .io_in2_im(BF_4_io_in2_im),
    .io_out1_re(BF_4_io_out1_re),
    .io_out1_im(BF_4_io_out1_im),
    .io_out2_re(BF_4_io_out2_re),
    .io_out2_im(BF_4_io_out2_im)
  );
  complexMul complexMul_4 ( // @[R2MDC.scala 60:22:@1221.4]
    .io_in1_re(complexMul_4_io_in1_re),
    .io_in1_im(complexMul_4_io_in1_im),
    .io_in2_re(complexMul_4_io_in2_re),
    .io_in2_im(complexMul_4_io_in2_im),
    .io_out_re(complexMul_4_io_out_re),
    .io_out_im(complexMul_4_io_out_im)
  );
  Switch Switch_4 ( // @[R2MDC.scala 80:22:@1234.4]
    .io_in1_re(Switch_4_io_in1_re),
    .io_in1_im(Switch_4_io_in1_im),
    .io_in2_re(Switch_4_io_in2_re),
    .io_in2_im(Switch_4_io_in2_im),
    .io_sel(Switch_4_io_sel),
    .io_out1_re(Switch_4_io_out1_re),
    .io_out1_im(Switch_4_io_out1_im),
    .io_out2_re(Switch_4_io_out2_re),
    .io_out2_im(Switch_4_io_out2_im)
  );
  BF BF_5 ( // @[R2MDC.scala 33:22:@1251.4]
    .io_in1_re(BF_5_io_in1_re),
    .io_in1_im(BF_5_io_in1_im),
    .io_in2_re(BF_5_io_in2_re),
    .io_in2_im(BF_5_io_in2_im),
    .io_out1_re(BF_5_io_out1_re),
    .io_out1_im(BF_5_io_out1_im),
    .io_out2_re(BF_5_io_out2_re),
    .io_out2_im(BF_5_io_out2_im)
  );
  assign _T_18 = cnt + 6'h1; // @[R2MDC.scala 122:16:@342.6]
  assign _T_19 = _T_18[5:0]; // @[R2MDC.scala 122:16:@343.6]
  assign _GEN_0 = io_din_valid ? _T_19 : cnt; // @[R2MDC.scala 121:21:@341.4]
  assign _T_239 = cnt[4:0]; // @[R2MDC.scala 131:23:@659.4]
  assign _GEN_66 = 5'h1 == _T_239 ? $signed(10'shff) : $signed(10'sh100); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_67 = 5'h2 == _T_239 ? $signed(10'shfb) : $signed(_GEN_66); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_68 = 5'h3 == _T_239 ? $signed(10'shf5) : $signed(_GEN_67); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_69 = 5'h4 == _T_239 ? $signed(10'shed) : $signed(_GEN_68); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_70 = 5'h5 == _T_239 ? $signed(10'she2) : $signed(_GEN_69); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_71 = 5'h6 == _T_239 ? $signed(10'shd5) : $signed(_GEN_70); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_72 = 5'h7 == _T_239 ? $signed(10'shc6) : $signed(_GEN_71); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_73 = 5'h8 == _T_239 ? $signed(10'shb5) : $signed(_GEN_72); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_74 = 5'h9 == _T_239 ? $signed(10'sha2) : $signed(_GEN_73); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_75 = 5'ha == _T_239 ? $signed(10'sh8e) : $signed(_GEN_74); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_76 = 5'hb == _T_239 ? $signed(10'sh79) : $signed(_GEN_75); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_77 = 5'hc == _T_239 ? $signed(10'sh62) : $signed(_GEN_76); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_78 = 5'hd == _T_239 ? $signed(10'sh4a) : $signed(_GEN_77); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_79 = 5'he == _T_239 ? $signed(10'sh32) : $signed(_GEN_78); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_80 = 5'hf == _T_239 ? $signed(10'sh19) : $signed(_GEN_79); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_81 = 5'h10 == _T_239 ? $signed(10'sh0) : $signed(_GEN_80); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_82 = 5'h11 == _T_239 ? $signed(-10'sh19) : $signed(_GEN_81); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_83 = 5'h12 == _T_239 ? $signed(-10'sh32) : $signed(_GEN_82); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_84 = 5'h13 == _T_239 ? $signed(-10'sh4a) : $signed(_GEN_83); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_85 = 5'h14 == _T_239 ? $signed(-10'sh62) : $signed(_GEN_84); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_86 = 5'h15 == _T_239 ? $signed(-10'sh79) : $signed(_GEN_85); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_87 = 5'h16 == _T_239 ? $signed(-10'sh8e) : $signed(_GEN_86); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_88 = 5'h17 == _T_239 ? $signed(-10'sha2) : $signed(_GEN_87); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_89 = 5'h18 == _T_239 ? $signed(-10'shb5) : $signed(_GEN_88); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_90 = 5'h19 == _T_239 ? $signed(-10'shc6) : $signed(_GEN_89); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_91 = 5'h1a == _T_239 ? $signed(-10'shd5) : $signed(_GEN_90); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_92 = 5'h1b == _T_239 ? $signed(-10'she2) : $signed(_GEN_91); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_93 = 5'h1c == _T_239 ? $signed(-10'shed) : $signed(_GEN_92); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_94 = 5'h1d == _T_239 ? $signed(-10'shf5) : $signed(_GEN_93); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_95 = 5'h1e == _T_239 ? $signed(-10'shfb) : $signed(_GEN_94); // @[R2MDC.scala 115:12:@694.4]
  assign _GEN_98 = 5'h1 == _T_239 ? $signed(-10'sh19) : $signed(10'sh0); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_99 = 5'h2 == _T_239 ? $signed(-10'sh32) : $signed(_GEN_98); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_100 = 5'h3 == _T_239 ? $signed(-10'sh4a) : $signed(_GEN_99); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_101 = 5'h4 == _T_239 ? $signed(-10'sh62) : $signed(_GEN_100); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_102 = 5'h5 == _T_239 ? $signed(-10'sh79) : $signed(_GEN_101); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_103 = 5'h6 == _T_239 ? $signed(-10'sh8e) : $signed(_GEN_102); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_104 = 5'h7 == _T_239 ? $signed(-10'sha2) : $signed(_GEN_103); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_105 = 5'h8 == _T_239 ? $signed(-10'shb5) : $signed(_GEN_104); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_106 = 5'h9 == _T_239 ? $signed(-10'shc6) : $signed(_GEN_105); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_107 = 5'ha == _T_239 ? $signed(-10'shd5) : $signed(_GEN_106); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_108 = 5'hb == _T_239 ? $signed(-10'she2) : $signed(_GEN_107); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_109 = 5'hc == _T_239 ? $signed(-10'shed) : $signed(_GEN_108); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_110 = 5'hd == _T_239 ? $signed(-10'shf5) : $signed(_GEN_109); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_111 = 5'he == _T_239 ? $signed(-10'shfb) : $signed(_GEN_110); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_112 = 5'hf == _T_239 ? $signed(-10'shff) : $signed(_GEN_111); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_113 = 5'h10 == _T_239 ? $signed(-10'sh100) : $signed(_GEN_112); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_114 = 5'h11 == _T_239 ? $signed(-10'shff) : $signed(_GEN_113); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_115 = 5'h12 == _T_239 ? $signed(-10'shfb) : $signed(_GEN_114); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_116 = 5'h13 == _T_239 ? $signed(-10'shf5) : $signed(_GEN_115); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_117 = 5'h14 == _T_239 ? $signed(-10'shed) : $signed(_GEN_116); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_118 = 5'h15 == _T_239 ? $signed(-10'she2) : $signed(_GEN_117); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_119 = 5'h16 == _T_239 ? $signed(-10'shd5) : $signed(_GEN_118); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_120 = 5'h17 == _T_239 ? $signed(-10'shc6) : $signed(_GEN_119); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_121 = 5'h18 == _T_239 ? $signed(-10'shb5) : $signed(_GEN_120); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_122 = 5'h19 == _T_239 ? $signed(-10'sha2) : $signed(_GEN_121); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_123 = 5'h1a == _T_239 ? $signed(-10'sh8e) : $signed(_GEN_122); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_124 = 5'h1b == _T_239 ? $signed(-10'sh79) : $signed(_GEN_123); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_125 = 5'h1c == _T_239 ? $signed(-10'sh62) : $signed(_GEN_124); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_126 = 5'h1d == _T_239 ? $signed(-10'sh4a) : $signed(_GEN_125); // @[R2MDC.scala 116:12:@728.4]
  assign _GEN_127 = 5'h1e == _T_239 ? $signed(-10'sh32) : $signed(_GEN_126); // @[R2MDC.scala 116:12:@728.4]
  assign _T_451 = cnt[3:0]; // @[R2MDC.scala 144:23:@916.4]
  assign _GEN_194 = 4'h1 == _T_451 ? $signed(10'shfb) : $signed(10'sh100); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_195 = 4'h2 == _T_451 ? $signed(10'shed) : $signed(_GEN_194); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_196 = 4'h3 == _T_451 ? $signed(10'shd5) : $signed(_GEN_195); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_197 = 4'h4 == _T_451 ? $signed(10'shb5) : $signed(_GEN_196); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_198 = 4'h5 == _T_451 ? $signed(10'sh8e) : $signed(_GEN_197); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_199 = 4'h6 == _T_451 ? $signed(10'sh62) : $signed(_GEN_198); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_200 = 4'h7 == _T_451 ? $signed(10'sh32) : $signed(_GEN_199); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_201 = 4'h8 == _T_451 ? $signed(10'sh0) : $signed(_GEN_200); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_202 = 4'h9 == _T_451 ? $signed(-10'sh32) : $signed(_GEN_201); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_203 = 4'ha == _T_451 ? $signed(-10'sh62) : $signed(_GEN_202); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_204 = 4'hb == _T_451 ? $signed(-10'sh8e) : $signed(_GEN_203); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_205 = 4'hc == _T_451 ? $signed(-10'shb5) : $signed(_GEN_204); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_206 = 4'hd == _T_451 ? $signed(-10'shd5) : $signed(_GEN_205); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_207 = 4'he == _T_451 ? $signed(-10'shed) : $signed(_GEN_206); // @[R2MDC.scala 115:12:@935.4]
  assign _GEN_210 = 4'h1 == _T_451 ? $signed(-10'sh32) : $signed(10'sh0); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_211 = 4'h2 == _T_451 ? $signed(-10'sh62) : $signed(_GEN_210); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_212 = 4'h3 == _T_451 ? $signed(-10'sh8e) : $signed(_GEN_211); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_213 = 4'h4 == _T_451 ? $signed(-10'shb5) : $signed(_GEN_212); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_214 = 4'h5 == _T_451 ? $signed(-10'shd5) : $signed(_GEN_213); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_215 = 4'h6 == _T_451 ? $signed(-10'shed) : $signed(_GEN_214); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_216 = 4'h7 == _T_451 ? $signed(-10'shfb) : $signed(_GEN_215); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_217 = 4'h8 == _T_451 ? $signed(-10'sh100) : $signed(_GEN_216); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_218 = 4'h9 == _T_451 ? $signed(-10'shfb) : $signed(_GEN_217); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_219 = 4'ha == _T_451 ? $signed(-10'shed) : $signed(_GEN_218); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_220 = 4'hb == _T_451 ? $signed(-10'shd5) : $signed(_GEN_219); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_221 = 4'hc == _T_451 ? $signed(-10'shb5) : $signed(_GEN_220); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_222 = 4'hd == _T_451 ? $signed(-10'sh8e) : $signed(_GEN_221); // @[R2MDC.scala 116:12:@953.4]
  assign _GEN_223 = 4'he == _T_451 ? $signed(-10'sh62) : $signed(_GEN_222); // @[R2MDC.scala 116:12:@953.4]
  assign _T_567 = cnt[2:0]; // @[R2MDC.scala 144:23:@1061.4]
  assign _GEN_258 = 3'h1 == _T_567 ? $signed(10'shed) : $signed(10'sh100); // @[R2MDC.scala 115:12:@1072.4]
  assign _GEN_259 = 3'h2 == _T_567 ? $signed(10'shb5) : $signed(_GEN_258); // @[R2MDC.scala 115:12:@1072.4]
  assign _GEN_260 = 3'h3 == _T_567 ? $signed(10'sh62) : $signed(_GEN_259); // @[R2MDC.scala 115:12:@1072.4]
  assign _GEN_261 = 3'h4 == _T_567 ? $signed(10'sh0) : $signed(_GEN_260); // @[R2MDC.scala 115:12:@1072.4]
  assign _GEN_262 = 3'h5 == _T_567 ? $signed(-10'sh62) : $signed(_GEN_261); // @[R2MDC.scala 115:12:@1072.4]
  assign _GEN_263 = 3'h6 == _T_567 ? $signed(-10'shb5) : $signed(_GEN_262); // @[R2MDC.scala 115:12:@1072.4]
  assign _GEN_266 = 3'h1 == _T_567 ? $signed(-10'sh62) : $signed(10'sh0); // @[R2MDC.scala 116:12:@1082.4]
  assign _GEN_267 = 3'h2 == _T_567 ? $signed(-10'shb5) : $signed(_GEN_266); // @[R2MDC.scala 116:12:@1082.4]
  assign _GEN_268 = 3'h3 == _T_567 ? $signed(-10'shed) : $signed(_GEN_267); // @[R2MDC.scala 116:12:@1082.4]
  assign _GEN_269 = 3'h4 == _T_567 ? $signed(-10'sh100) : $signed(_GEN_268); // @[R2MDC.scala 116:12:@1082.4]
  assign _GEN_270 = 3'h5 == _T_567 ? $signed(-10'shed) : $signed(_GEN_269); // @[R2MDC.scala 116:12:@1082.4]
  assign _GEN_271 = 3'h6 == _T_567 ? $signed(-10'shb5) : $signed(_GEN_270); // @[R2MDC.scala 116:12:@1082.4]
  assign _T_635 = cnt[1:0]; // @[R2MDC.scala 144:23:@1150.4]
  assign _GEN_290 = 2'h1 == _T_635 ? $signed(10'shb5) : $signed(10'sh100); // @[R2MDC.scala 115:12:@1157.4]
  assign _GEN_291 = 2'h2 == _T_635 ? $signed(10'sh0) : $signed(_GEN_290); // @[R2MDC.scala 115:12:@1157.4]
  assign _GEN_294 = 2'h1 == _T_635 ? $signed(-10'shb5) : $signed(10'sh0); // @[R2MDC.scala 116:12:@1163.4]
  assign _GEN_295 = 2'h2 == _T_635 ? $signed(-10'sh100) : $signed(_GEN_294); // @[R2MDC.scala 116:12:@1163.4]
  assign _T_679 = cnt[0]; // @[R2MDC.scala 144:23:@1211.4]
  assign io_dOut1_re = _T_712_re; // @[R2MDC.scala 161:12:@1266.4]
  assign io_dOut1_im = _T_712_im; // @[R2MDC.scala 161:12:@1265.4]
  assign io_dOut2_re = _T_714_re; // @[R2MDC.scala 162:12:@1271.4]
  assign io_dOut2_im = _T_714_im; // @[R2MDC.scala 162:12:@1270.4]
  assign io_dout_valid = _T_843; // @[R2MDC.scala 163:17:@1528.4]
  assign BF_io_in1_re = _T_238_re; // @[R2MDC.scala 34:17:@656.4]
  assign BF_io_in1_im = _T_238_im; // @[R2MDC.scala 34:17:@655.4]
  assign BF_io_in2_re = io_dIn_re; // @[R2MDC.scala 35:17:@658.4]
  assign BF_io_in2_im = io_dIn_im; // @[R2MDC.scala 35:17:@657.4]
  assign complexMul_io_in1_re = BF_io_out2_re; // @[R2MDC.scala 61:17:@733.4]
  assign complexMul_io_in1_im = BF_io_out2_im; // @[R2MDC.scala 61:17:@732.4]
  assign complexMul_io_in2_re = 5'h1f == _T_239 ? $signed(-10'shff) : $signed(_GEN_95); // @[R2MDC.scala 62:17:@735.4]
  assign complexMul_io_in2_im = 5'h1f == _T_239 ? $signed(-10'sh19) : $signed(_GEN_127); // @[R2MDC.scala 62:17:@734.4]
  assign Switch_io_in1_re = BF_io_out1_re; // @[R2MDC.scala 81:17:@821.4]
  assign Switch_io_in1_im = BF_io_out1_im; // @[R2MDC.scala 81:17:@820.4]
  assign Switch_io_in2_re = _T_416_re; // @[R2MDC.scala 82:17:@823.4]
  assign Switch_io_in2_im = _T_416_im; // @[R2MDC.scala 82:17:@822.4]
  assign Switch_io_sel = cnt[4]; // @[R2MDC.scala 83:17:@824.4]
  assign BF_1_io_in1_re = _T_450_re; // @[R2MDC.scala 34:17:@913.4]
  assign BF_1_io_in1_im = _T_450_im; // @[R2MDC.scala 34:17:@912.4]
  assign BF_1_io_in2_re = Switch_io_out2_re; // @[R2MDC.scala 35:17:@915.4]
  assign BF_1_io_in2_im = Switch_io_out2_im; // @[R2MDC.scala 35:17:@914.4]
  assign complexMul_1_io_in1_re = BF_1_io_out2_re; // @[R2MDC.scala 61:17:@958.4]
  assign complexMul_1_io_in1_im = BF_1_io_out2_im; // @[R2MDC.scala 61:17:@957.4]
  assign complexMul_1_io_in2_re = 4'hf == _T_451 ? $signed(-10'shfb) : $signed(_GEN_207); // @[R2MDC.scala 62:17:@960.4]
  assign complexMul_1_io_in2_im = 4'hf == _T_451 ? $signed(-10'sh32) : $signed(_GEN_223); // @[R2MDC.scala 62:17:@959.4]
  assign Switch_1_io_in1_re = BF_1_io_out1_re; // @[R2MDC.scala 81:17:@1006.4]
  assign Switch_1_io_in1_im = BF_1_io_out1_im; // @[R2MDC.scala 81:17:@1005.4]
  assign Switch_1_io_in2_re = _T_548_re; // @[R2MDC.scala 82:17:@1008.4]
  assign Switch_1_io_in2_im = _T_548_im; // @[R2MDC.scala 82:17:@1007.4]
  assign Switch_1_io_sel = cnt[3]; // @[R2MDC.scala 83:17:@1009.4]
  assign BF_2_io_in1_re = _T_566_re; // @[R2MDC.scala 34:17:@1058.4]
  assign BF_2_io_in1_im = _T_566_im; // @[R2MDC.scala 34:17:@1057.4]
  assign BF_2_io_in2_re = Switch_1_io_out2_re; // @[R2MDC.scala 35:17:@1060.4]
  assign BF_2_io_in2_im = Switch_1_io_out2_im; // @[R2MDC.scala 35:17:@1059.4]
  assign complexMul_2_io_in1_re = BF_2_io_out2_re; // @[R2MDC.scala 61:17:@1087.4]
  assign complexMul_2_io_in1_im = BF_2_io_out2_im; // @[R2MDC.scala 61:17:@1086.4]
  assign complexMul_2_io_in2_re = 3'h7 == _T_567 ? $signed(-10'shed) : $signed(_GEN_263); // @[R2MDC.scala 62:17:@1089.4]
  assign complexMul_2_io_in2_im = 3'h7 == _T_567 ? $signed(-10'sh62) : $signed(_GEN_271); // @[R2MDC.scala 62:17:@1088.4]
  assign Switch_2_io_in1_re = BF_2_io_out1_re; // @[R2MDC.scala 81:17:@1115.4]
  assign Switch_2_io_in1_im = BF_2_io_out1_im; // @[R2MDC.scala 81:17:@1114.4]
  assign Switch_2_io_in2_re = _T_624_re; // @[R2MDC.scala 82:17:@1117.4]
  assign Switch_2_io_in2_im = _T_624_im; // @[R2MDC.scala 82:17:@1116.4]
  assign Switch_2_io_sel = cnt[2]; // @[R2MDC.scala 83:17:@1118.4]
  assign BF_3_io_in1_re = _T_634_re; // @[R2MDC.scala 34:17:@1147.4]
  assign BF_3_io_in1_im = _T_634_im; // @[R2MDC.scala 34:17:@1146.4]
  assign BF_3_io_in2_re = Switch_2_io_out2_re; // @[R2MDC.scala 35:17:@1149.4]
  assign BF_3_io_in2_im = Switch_2_io_out2_im; // @[R2MDC.scala 35:17:@1148.4]
  assign complexMul_3_io_in1_re = BF_3_io_out2_re; // @[R2MDC.scala 61:17:@1168.4]
  assign complexMul_3_io_in1_im = BF_3_io_out2_im; // @[R2MDC.scala 61:17:@1167.4]
  assign complexMul_3_io_in2_re = 2'h3 == _T_635 ? $signed(-10'shb5) : $signed(_GEN_291); // @[R2MDC.scala 62:17:@1170.4]
  assign complexMul_3_io_in2_im = 2'h3 == _T_635 ? $signed(-10'shb5) : $signed(_GEN_295); // @[R2MDC.scala 62:17:@1169.4]
  assign Switch_3_io_in1_re = BF_3_io_out1_re; // @[R2MDC.scala 81:17:@1186.4]
  assign Switch_3_io_in1_im = BF_3_io_out1_im; // @[R2MDC.scala 81:17:@1185.4]
  assign Switch_3_io_in2_re = _T_672_re; // @[R2MDC.scala 82:17:@1188.4]
  assign Switch_3_io_in2_im = _T_672_im; // @[R2MDC.scala 82:17:@1187.4]
  assign Switch_3_io_sel = cnt[1]; // @[R2MDC.scala 83:17:@1189.4]
  assign BF_4_io_in1_re = _T_678_re; // @[R2MDC.scala 34:17:@1208.4]
  assign BF_4_io_in1_im = _T_678_im; // @[R2MDC.scala 34:17:@1207.4]
  assign BF_4_io_in2_re = Switch_3_io_out2_re; // @[R2MDC.scala 35:17:@1210.4]
  assign BF_4_io_in2_im = Switch_3_io_out2_im; // @[R2MDC.scala 35:17:@1209.4]
  assign complexMul_4_io_in1_re = BF_4_io_out2_re; // @[R2MDC.scala 61:17:@1225.4]
  assign complexMul_4_io_in1_im = BF_4_io_out2_im; // @[R2MDC.scala 61:17:@1224.4]
  assign complexMul_4_io_in2_re = _T_679 ? $signed(10'sh0) : $signed(10'sh100); // @[R2MDC.scala 62:17:@1227.4]
  assign complexMul_4_io_in2_im = _T_679 ? $signed(-10'sh100) : $signed(10'sh0); // @[R2MDC.scala 62:17:@1226.4]
  assign Switch_4_io_in1_re = BF_4_io_out1_re; // @[R2MDC.scala 81:17:@1238.4]
  assign Switch_4_io_in1_im = BF_4_io_out1_im; // @[R2MDC.scala 81:17:@1237.4]
  assign Switch_4_io_in2_re = _T_706_re; // @[R2MDC.scala 82:17:@1240.4]
  assign Switch_4_io_in2_im = _T_706_im; // @[R2MDC.scala 82:17:@1239.4]
  assign Switch_4_io_sel = cnt[0]; // @[R2MDC.scala 83:17:@1241.4]
  assign BF_5_io_in1_re = _T_710_re; // @[R2MDC.scala 34:17:@1255.4]
  assign BF_5_io_in1_im = _T_710_im; // @[R2MDC.scala 34:17:@1254.4]
  assign BF_5_io_in2_re = Switch_4_io_out2_re; // @[R2MDC.scala 35:17:@1257.4]
  assign BF_5_io_in2_im = Switch_4_io_out2_im; // @[R2MDC.scala 35:17:@1256.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_176_re = _RAND_1[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_176_im = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_178_re = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_178_im = _RAND_4[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_180_re = _RAND_5[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_180_im = _RAND_6[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_182_re = _RAND_7[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_182_im = _RAND_8[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_184_re = _RAND_9[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_184_im = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_186_re = _RAND_11[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_186_im = _RAND_12[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_188_re = _RAND_13[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_188_im = _RAND_14[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_190_re = _RAND_15[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_190_im = _RAND_16[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_192_re = _RAND_17[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_192_im = _RAND_18[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_194_re = _RAND_19[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_194_im = _RAND_20[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_196_re = _RAND_21[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_196_im = _RAND_22[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_198_re = _RAND_23[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_198_im = _RAND_24[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_200_re = _RAND_25[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_200_im = _RAND_26[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_202_re = _RAND_27[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_202_im = _RAND_28[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_204_re = _RAND_29[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_204_im = _RAND_30[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_206_re = _RAND_31[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_206_im = _RAND_32[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_208_re = _RAND_33[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_208_im = _RAND_34[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_210_re = _RAND_35[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_210_im = _RAND_36[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_212_re = _RAND_37[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_212_im = _RAND_38[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_214_re = _RAND_39[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_214_im = _RAND_40[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_216_re = _RAND_41[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_216_im = _RAND_42[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_218_re = _RAND_43[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_218_im = _RAND_44[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_220_re = _RAND_45[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_220_im = _RAND_46[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_222_re = _RAND_47[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_222_im = _RAND_48[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_224_re = _RAND_49[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_224_im = _RAND_50[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_226_re = _RAND_51[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_226_im = _RAND_52[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_228_re = _RAND_53[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_228_im = _RAND_54[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_230_re = _RAND_55[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_230_im = _RAND_56[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_232_re = _RAND_57[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_232_im = _RAND_58[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_234_re = _RAND_59[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_234_im = _RAND_60[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_236_re = _RAND_61[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_236_im = _RAND_62[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_238_re = _RAND_63[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_238_im = _RAND_64[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_386_re = _RAND_65[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_386_im = _RAND_66[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_388_re = _RAND_67[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_388_im = _RAND_68[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_390_re = _RAND_69[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_390_im = _RAND_70[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_392_re = _RAND_71[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_392_im = _RAND_72[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_394_re = _RAND_73[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_394_im = _RAND_74[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_396_re = _RAND_75[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_396_im = _RAND_76[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_398_re = _RAND_77[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_398_im = _RAND_78[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_400_re = _RAND_79[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_400_im = _RAND_80[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_402_re = _RAND_81[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_402_im = _RAND_82[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_404_re = _RAND_83[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_404_im = _RAND_84[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_406_re = _RAND_85[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_406_im = _RAND_86[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_408_re = _RAND_87[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_408_im = _RAND_88[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_410_re = _RAND_89[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_410_im = _RAND_90[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_412_re = _RAND_91[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_412_im = _RAND_92[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_414_re = _RAND_93[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_414_im = _RAND_94[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_416_re = _RAND_95[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_416_im = _RAND_96[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_420_re = _RAND_97[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_420_im = _RAND_98[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_422_re = _RAND_99[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_422_im = _RAND_100[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_424_re = _RAND_101[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_424_im = _RAND_102[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_426_re = _RAND_103[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_426_im = _RAND_104[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_428_re = _RAND_105[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_428_im = _RAND_106[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_430_re = _RAND_107[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_430_im = _RAND_108[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_432_re = _RAND_109[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_432_im = _RAND_110[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_434_re = _RAND_111[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_434_im = _RAND_112[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_436_re = _RAND_113[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_436_im = _RAND_114[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_438_re = _RAND_115[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_438_im = _RAND_116[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_440_re = _RAND_117[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_440_im = _RAND_118[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_442_re = _RAND_119[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_442_im = _RAND_120[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_444_re = _RAND_121[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_444_im = _RAND_122[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_446_re = _RAND_123[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_446_im = _RAND_124[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_448_re = _RAND_125[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_448_im = _RAND_126[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_450_re = _RAND_127[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_450_im = _RAND_128[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_534_re = _RAND_129[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_534_im = _RAND_130[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_536_re = _RAND_131[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_536_im = _RAND_132[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_538_re = _RAND_133[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_538_im = _RAND_134[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_540_re = _RAND_135[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_540_im = _RAND_136[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_542_re = _RAND_137[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_542_im = _RAND_138[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_544_re = _RAND_139[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_544_im = _RAND_140[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_546_re = _RAND_141[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_546_im = _RAND_142[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_548_re = _RAND_143[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_548_im = _RAND_144[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_552_re = _RAND_145[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_552_im = _RAND_146[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_554_re = _RAND_147[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_554_im = _RAND_148[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_556_re = _RAND_149[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_556_im = _RAND_150[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_558_re = _RAND_151[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_558_im = _RAND_152[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_560_re = _RAND_153[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_560_im = _RAND_154[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_562_re = _RAND_155[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_562_im = _RAND_156[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_564_re = _RAND_157[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_564_im = _RAND_158[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_566_re = _RAND_159[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_566_im = _RAND_160[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_618_re = _RAND_161[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_618_im = _RAND_162[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_620_re = _RAND_163[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_620_im = _RAND_164[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_622_re = _RAND_165[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_622_im = _RAND_166[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_624_re = _RAND_167[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_624_im = _RAND_168[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_628_re = _RAND_169[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_628_im = _RAND_170[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_630_re = _RAND_171[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_630_im = _RAND_172[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_632_re = _RAND_173[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_632_im = _RAND_174[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_634_re = _RAND_175[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_634_im = _RAND_176[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_670_re = _RAND_177[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_670_im = _RAND_178[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_672_re = _RAND_179[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_672_im = _RAND_180[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_676_re = _RAND_181[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_676_im = _RAND_182[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_678_re = _RAND_183[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_678_im = _RAND_184[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_706_re = _RAND_185[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_706_im = _RAND_186[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_710_re = _RAND_187[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_710_im = _RAND_188[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_712_re = _RAND_189[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_712_im = _RAND_190[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_714_re = _RAND_191[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_714_im = _RAND_192[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_717 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_719 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_721 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_723 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_725 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_727 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_729 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_731 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_733 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_735 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_737 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_739 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_741 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_743 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_745 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_747 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_749 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_751 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_753 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_755 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_757 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_759 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_761 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_763 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_765 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_767 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_769 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_771 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_773 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_775 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_777 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_779 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_781 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_783 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_785 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_787 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_789 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_791 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_793 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_795 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_797 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_799 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_801 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_803 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_805 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_807 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_809 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_811 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_813 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_815 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_817 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_819 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_821 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_823 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_825 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_827 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_829 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_831 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_833 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_835 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_837 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_839 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_841 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_843 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 6'h0;
    end else begin
      if (io_din_valid) begin
        cnt <= _T_19;
      end
    end
    _T_176_re <= io_dIn_re;
    _T_176_im <= io_dIn_im;
    _T_178_re <= _T_176_re;
    _T_178_im <= _T_176_im;
    _T_180_re <= _T_178_re;
    _T_180_im <= _T_178_im;
    _T_182_re <= _T_180_re;
    _T_182_im <= _T_180_im;
    _T_184_re <= _T_182_re;
    _T_184_im <= _T_182_im;
    _T_186_re <= _T_184_re;
    _T_186_im <= _T_184_im;
    _T_188_re <= _T_186_re;
    _T_188_im <= _T_186_im;
    _T_190_re <= _T_188_re;
    _T_190_im <= _T_188_im;
    _T_192_re <= _T_190_re;
    _T_192_im <= _T_190_im;
    _T_194_re <= _T_192_re;
    _T_194_im <= _T_192_im;
    _T_196_re <= _T_194_re;
    _T_196_im <= _T_194_im;
    _T_198_re <= _T_196_re;
    _T_198_im <= _T_196_im;
    _T_200_re <= _T_198_re;
    _T_200_im <= _T_198_im;
    _T_202_re <= _T_200_re;
    _T_202_im <= _T_200_im;
    _T_204_re <= _T_202_re;
    _T_204_im <= _T_202_im;
    _T_206_re <= _T_204_re;
    _T_206_im <= _T_204_im;
    _T_208_re <= _T_206_re;
    _T_208_im <= _T_206_im;
    _T_210_re <= _T_208_re;
    _T_210_im <= _T_208_im;
    _T_212_re <= _T_210_re;
    _T_212_im <= _T_210_im;
    _T_214_re <= _T_212_re;
    _T_214_im <= _T_212_im;
    _T_216_re <= _T_214_re;
    _T_216_im <= _T_214_im;
    _T_218_re <= _T_216_re;
    _T_218_im <= _T_216_im;
    _T_220_re <= _T_218_re;
    _T_220_im <= _T_218_im;
    _T_222_re <= _T_220_re;
    _T_222_im <= _T_220_im;
    _T_224_re <= _T_222_re;
    _T_224_im <= _T_222_im;
    _T_226_re <= _T_224_re;
    _T_226_im <= _T_224_im;
    _T_228_re <= _T_226_re;
    _T_228_im <= _T_226_im;
    _T_230_re <= _T_228_re;
    _T_230_im <= _T_228_im;
    _T_232_re <= _T_230_re;
    _T_232_im <= _T_230_im;
    _T_234_re <= _T_232_re;
    _T_234_im <= _T_232_im;
    _T_236_re <= _T_234_re;
    _T_236_im <= _T_234_im;
    _T_238_re <= _T_236_re;
    _T_238_im <= _T_236_im;
    _T_386_re <= complexMul_io_out_re;
    _T_386_im <= complexMul_io_out_im;
    _T_388_re <= _T_386_re;
    _T_388_im <= _T_386_im;
    _T_390_re <= _T_388_re;
    _T_390_im <= _T_388_im;
    _T_392_re <= _T_390_re;
    _T_392_im <= _T_390_im;
    _T_394_re <= _T_392_re;
    _T_394_im <= _T_392_im;
    _T_396_re <= _T_394_re;
    _T_396_im <= _T_394_im;
    _T_398_re <= _T_396_re;
    _T_398_im <= _T_396_im;
    _T_400_re <= _T_398_re;
    _T_400_im <= _T_398_im;
    _T_402_re <= _T_400_re;
    _T_402_im <= _T_400_im;
    _T_404_re <= _T_402_re;
    _T_404_im <= _T_402_im;
    _T_406_re <= _T_404_re;
    _T_406_im <= _T_404_im;
    _T_408_re <= _T_406_re;
    _T_408_im <= _T_406_im;
    _T_410_re <= _T_408_re;
    _T_410_im <= _T_408_im;
    _T_412_re <= _T_410_re;
    _T_412_im <= _T_410_im;
    _T_414_re <= _T_412_re;
    _T_414_im <= _T_412_im;
    _T_416_re <= _T_414_re;
    _T_416_im <= _T_414_im;
    _T_420_re <= Switch_io_out1_re;
    _T_420_im <= Switch_io_out1_im;
    _T_422_re <= _T_420_re;
    _T_422_im <= _T_420_im;
    _T_424_re <= _T_422_re;
    _T_424_im <= _T_422_im;
    _T_426_re <= _T_424_re;
    _T_426_im <= _T_424_im;
    _T_428_re <= _T_426_re;
    _T_428_im <= _T_426_im;
    _T_430_re <= _T_428_re;
    _T_430_im <= _T_428_im;
    _T_432_re <= _T_430_re;
    _T_432_im <= _T_430_im;
    _T_434_re <= _T_432_re;
    _T_434_im <= _T_432_im;
    _T_436_re <= _T_434_re;
    _T_436_im <= _T_434_im;
    _T_438_re <= _T_436_re;
    _T_438_im <= _T_436_im;
    _T_440_re <= _T_438_re;
    _T_440_im <= _T_438_im;
    _T_442_re <= _T_440_re;
    _T_442_im <= _T_440_im;
    _T_444_re <= _T_442_re;
    _T_444_im <= _T_442_im;
    _T_446_re <= _T_444_re;
    _T_446_im <= _T_444_im;
    _T_448_re <= _T_446_re;
    _T_448_im <= _T_446_im;
    _T_450_re <= _T_448_re;
    _T_450_im <= _T_448_im;
    _T_534_re <= complexMul_1_io_out_re;
    _T_534_im <= complexMul_1_io_out_im;
    _T_536_re <= _T_534_re;
    _T_536_im <= _T_534_im;
    _T_538_re <= _T_536_re;
    _T_538_im <= _T_536_im;
    _T_540_re <= _T_538_re;
    _T_540_im <= _T_538_im;
    _T_542_re <= _T_540_re;
    _T_542_im <= _T_540_im;
    _T_544_re <= _T_542_re;
    _T_544_im <= _T_542_im;
    _T_546_re <= _T_544_re;
    _T_546_im <= _T_544_im;
    _T_548_re <= _T_546_re;
    _T_548_im <= _T_546_im;
    _T_552_re <= Switch_1_io_out1_re;
    _T_552_im <= Switch_1_io_out1_im;
    _T_554_re <= _T_552_re;
    _T_554_im <= _T_552_im;
    _T_556_re <= _T_554_re;
    _T_556_im <= _T_554_im;
    _T_558_re <= _T_556_re;
    _T_558_im <= _T_556_im;
    _T_560_re <= _T_558_re;
    _T_560_im <= _T_558_im;
    _T_562_re <= _T_560_re;
    _T_562_im <= _T_560_im;
    _T_564_re <= _T_562_re;
    _T_564_im <= _T_562_im;
    _T_566_re <= _T_564_re;
    _T_566_im <= _T_564_im;
    _T_618_re <= complexMul_2_io_out_re;
    _T_618_im <= complexMul_2_io_out_im;
    _T_620_re <= _T_618_re;
    _T_620_im <= _T_618_im;
    _T_622_re <= _T_620_re;
    _T_622_im <= _T_620_im;
    _T_624_re <= _T_622_re;
    _T_624_im <= _T_622_im;
    _T_628_re <= Switch_2_io_out1_re;
    _T_628_im <= Switch_2_io_out1_im;
    _T_630_re <= _T_628_re;
    _T_630_im <= _T_628_im;
    _T_632_re <= _T_630_re;
    _T_632_im <= _T_630_im;
    _T_634_re <= _T_632_re;
    _T_634_im <= _T_632_im;
    _T_670_re <= complexMul_3_io_out_re;
    _T_670_im <= complexMul_3_io_out_im;
    _T_672_re <= _T_670_re;
    _T_672_im <= _T_670_im;
    _T_676_re <= Switch_3_io_out1_re;
    _T_676_im <= Switch_3_io_out1_im;
    _T_678_re <= _T_676_re;
    _T_678_im <= _T_676_im;
    _T_706_re <= complexMul_4_io_out_re;
    _T_706_im <= complexMul_4_io_out_im;
    _T_710_re <= Switch_4_io_out1_re;
    _T_710_im <= Switch_4_io_out1_im;
    _T_712_re <= BF_5_io_out1_re;
    _T_712_im <= BF_5_io_out1_im;
    _T_714_re <= BF_5_io_out2_re;
    _T_714_im <= BF_5_io_out2_im;
    _T_717 <= io_din_valid;
    _T_719 <= _T_717;
    _T_721 <= _T_719;
    _T_723 <= _T_721;
    _T_725 <= _T_723;
    _T_727 <= _T_725;
    _T_729 <= _T_727;
    _T_731 <= _T_729;
    _T_733 <= _T_731;
    _T_735 <= _T_733;
    _T_737 <= _T_735;
    _T_739 <= _T_737;
    _T_741 <= _T_739;
    _T_743 <= _T_741;
    _T_745 <= _T_743;
    _T_747 <= _T_745;
    _T_749 <= _T_747;
    _T_751 <= _T_749;
    _T_753 <= _T_751;
    _T_755 <= _T_753;
    _T_757 <= _T_755;
    _T_759 <= _T_757;
    _T_761 <= _T_759;
    _T_763 <= _T_761;
    _T_765 <= _T_763;
    _T_767 <= _T_765;
    _T_769 <= _T_767;
    _T_771 <= _T_769;
    _T_773 <= _T_771;
    _T_775 <= _T_773;
    _T_777 <= _T_775;
    _T_779 <= _T_777;
    _T_781 <= _T_779;
    _T_783 <= _T_781;
    _T_785 <= _T_783;
    _T_787 <= _T_785;
    _T_789 <= _T_787;
    _T_791 <= _T_789;
    _T_793 <= _T_791;
    _T_795 <= _T_793;
    _T_797 <= _T_795;
    _T_799 <= _T_797;
    _T_801 <= _T_799;
    _T_803 <= _T_801;
    _T_805 <= _T_803;
    _T_807 <= _T_805;
    _T_809 <= _T_807;
    _T_811 <= _T_809;
    _T_813 <= _T_811;
    _T_815 <= _T_813;
    _T_817 <= _T_815;
    _T_819 <= _T_817;
    _T_821 <= _T_819;
    _T_823 <= _T_821;
    _T_825 <= _T_823;
    _T_827 <= _T_825;
    _T_829 <= _T_827;
    _T_831 <= _T_829;
    _T_833 <= _T_831;
    _T_835 <= _T_833;
    _T_837 <= _T_835;
    _T_839 <= _T_837;
    _T_841 <= _T_839;
    _T_843 <= _T_841;
  end
endmodule
