module MR( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [27:0] io_a, // @[:@6.4]
  output [13:0] io_ar // @[:@6.4]
);
  wire [27:0] shift1; // @[MR.scala 26:21:@8.4]
  wire [28:0] _GEN_0; // @[MR.scala 27:31:@9.4]
  wire [28:0] _T_11; // @[MR.scala 27:31:@9.4]
  wire [29:0] _T_12; // @[MR.scala 27:21:@10.4]
  wire [28:0] _T_13; // @[MR.scala 27:21:@11.4]
  wire [30:0] _GEN_2; // @[MR.scala 27:49:@12.4]
  wire [30:0] _T_15; // @[MR.scala 27:49:@12.4]
  wire [30:0] _GEN_3; // @[MR.scala 27:39:@13.4]
  wire [31:0] _T_16; // @[MR.scala 27:39:@13.4]
  wire [30:0] _T_17; // @[MR.scala 27:39:@14.4]
  wire [34:0] _GEN_4; // @[MR.scala 27:67:@15.4]
  wire [34:0] _T_19; // @[MR.scala 27:67:@15.4]
  wire [34:0] _GEN_5; // @[MR.scala 27:57:@16.4]
  wire [35:0] _T_20; // @[MR.scala 27:57:@16.4]
  wire [34:0] _T_21; // @[MR.scala 27:57:@17.4]
  wire [34:0] _T_23; // @[MR.scala 27:85:@18.4]
  wire [35:0] _T_24; // @[MR.scala 27:75:@19.4]
  wire [34:0] _T_25; // @[MR.scala 27:75:@20.4]
  wire [42:0] _GEN_7; // @[MR.scala 28:13:@21.4]
  wire [42:0] _T_27; // @[MR.scala 28:13:@21.4]
  wire [42:0] _GEN_8; // @[MR.scala 27:93:@22.4]
  wire [43:0] _T_28; // @[MR.scala 27:93:@22.4]
  wire [42:0] _T_29; // @[MR.scala 27:93:@23.4]
  wire [42:0] _T_31; // @[MR.scala 28:31:@24.4]
  wire [43:0] _T_32; // @[MR.scala 28:21:@25.4]
  wire [42:0] _T_33; // @[MR.scala 28:21:@26.4]
  wire [42:0] _T_35; // @[MR.scala 28:50:@27.4]
  wire [43:0] _T_36; // @[MR.scala 28:40:@28.4]
  wire [42:0] _T_37; // @[MR.scala 28:40:@29.4]
  wire [42:0] _T_39; // @[MR.scala 28:69:@30.4]
  wire [43:0] _T_40; // @[MR.scala 28:59:@31.4]
  wire [42:0] mul1; // @[MR.scala 28:59:@32.4]
  wire [42:0] qGuess; // @[MR.scala 29:21:@33.4]
  wire [57:0] _GEN_12; // @[MR.scala 30:29:@34.4]
  wire [57:0] _T_43; // @[MR.scala 30:29:@34.4]
  wire [58:0] _T_44; // @[MR.scala 30:19:@35.4]
  wire [57:0] _T_45; // @[MR.scala 30:19:@36.4]
  wire [57:0] _T_47; // @[MR.scala 30:48:@37.4]
  wire [58:0] _T_48; // @[MR.scala 30:38:@38.4]
  wire [57:0] qM; // @[MR.scala 30:38:@39.4]
  wire [57:0] _GEN_15; // @[MR.scala 31:16:@40.4]
  wire [58:0] _T_49; // @[MR.scala 31:16:@40.4]
  wire [58:0] _T_50; // @[MR.scala 31:16:@41.4]
  wire [57:0] z; // @[MR.scala 31:16:@42.4]
  wire  _T_52; // @[MR.scala 32:18:@43.4]
  wire [58:0] _T_54; // @[MR.scala 32:45:@44.4]
  wire [58:0] _T_55; // @[MR.scala 32:45:@45.4]
  wire [57:0] _T_56; // @[MR.scala 32:45:@46.4]
  wire [57:0] _T_57; // @[MR.scala 32:15:@47.4]
  assign shift1 = io_a >> 4'hc; // @[MR.scala 26:21:@8.4]
  assign _GEN_0 = {{1'd0}, shift1}; // @[MR.scala 27:31:@9.4]
  assign _T_11 = _GEN_0 << 1'h1; // @[MR.scala 27:31:@9.4]
  assign _T_12 = _GEN_0 + _T_11; // @[MR.scala 27:21:@10.4]
  assign _T_13 = _T_12[28:0]; // @[MR.scala 27:21:@11.4]
  assign _GEN_2 = {{3'd0}, shift1}; // @[MR.scala 27:49:@12.4]
  assign _T_15 = _GEN_2 << 2'h2; // @[MR.scala 27:49:@12.4]
  assign _GEN_3 = {{2'd0}, _T_13}; // @[MR.scala 27:39:@13.4]
  assign _T_16 = _GEN_3 + _T_15; // @[MR.scala 27:39:@13.4]
  assign _T_17 = _T_16[30:0]; // @[MR.scala 27:39:@14.4]
  assign _GEN_4 = {{7'd0}, shift1}; // @[MR.scala 27:67:@15.4]
  assign _T_19 = _GEN_4 << 3'h5; // @[MR.scala 27:67:@15.4]
  assign _GEN_5 = {{4'd0}, _T_17}; // @[MR.scala 27:57:@16.4]
  assign _T_20 = _GEN_5 + _T_19; // @[MR.scala 27:57:@16.4]
  assign _T_21 = _T_20[34:0]; // @[MR.scala 27:57:@17.4]
  assign _T_23 = _GEN_4 << 3'h7; // @[MR.scala 27:85:@18.4]
  assign _T_24 = _T_21 + _T_23; // @[MR.scala 27:75:@19.4]
  assign _T_25 = _T_24[34:0]; // @[MR.scala 27:75:@20.4]
  assign _GEN_7 = {{15'd0}, shift1}; // @[MR.scala 28:13:@21.4]
  assign _T_27 = _GEN_7 << 4'h9; // @[MR.scala 28:13:@21.4]
  assign _GEN_8 = {{8'd0}, _T_25}; // @[MR.scala 27:93:@22.4]
  assign _T_28 = _GEN_8 + _T_27; // @[MR.scala 27:93:@22.4]
  assign _T_29 = _T_28[42:0]; // @[MR.scala 27:93:@23.4]
  assign _T_31 = _GEN_7 << 4'hb; // @[MR.scala 28:31:@24.4]
  assign _T_32 = _T_29 + _T_31; // @[MR.scala 28:21:@25.4]
  assign _T_33 = _T_32[42:0]; // @[MR.scala 28:21:@26.4]
  assign _T_35 = _GEN_7 << 4'hd; // @[MR.scala 28:50:@27.4]
  assign _T_36 = _T_33 + _T_35; // @[MR.scala 28:40:@28.4]
  assign _T_37 = _T_36[42:0]; // @[MR.scala 28:40:@29.4]
  assign _T_39 = _GEN_7 << 4'hf; // @[MR.scala 28:69:@30.4]
  assign _T_40 = _T_37 + _T_39; // @[MR.scala 28:59:@31.4]
  assign mul1 = _T_40[42:0]; // @[MR.scala 28:59:@32.4]
  assign qGuess = mul1 >> 5'h11; // @[MR.scala 29:21:@33.4]
  assign _GEN_12 = {{15'd0}, qGuess}; // @[MR.scala 30:29:@34.4]
  assign _T_43 = _GEN_12 << 4'hc; // @[MR.scala 30:29:@34.4]
  assign _T_44 = _GEN_12 + _T_43; // @[MR.scala 30:19:@35.4]
  assign _T_45 = _T_44[57:0]; // @[MR.scala 30:19:@36.4]
  assign _T_47 = _GEN_12 << 4'hd; // @[MR.scala 30:48:@37.4]
  assign _T_48 = _T_45 + _T_47; // @[MR.scala 30:38:@38.4]
  assign qM = _T_48[57:0]; // @[MR.scala 30:38:@39.4]
  assign _GEN_15 = {{30'd0}, io_a}; // @[MR.scala 31:16:@40.4]
  assign _T_49 = _GEN_15 - qM; // @[MR.scala 31:16:@40.4]
  assign _T_50 = $unsigned(_T_49); // @[MR.scala 31:16:@41.4]
  assign z = _T_50[57:0]; // @[MR.scala 31:16:@42.4]
  assign _T_52 = z < 58'h3001; // @[MR.scala 32:18:@43.4]
  assign _T_54 = z - 58'h3001; // @[MR.scala 32:45:@44.4]
  assign _T_55 = $unsigned(_T_54); // @[MR.scala 32:45:@45.4]
  assign _T_56 = _T_55[57:0]; // @[MR.scala 32:45:@46.4]
  assign _T_57 = _T_52 ? z : _T_56; // @[MR.scala 32:15:@47.4]
  assign io_ar = _T_57[13:0]; // @[MR.scala 32:9:@48.4]
endmodule
