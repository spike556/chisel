module OneBit( // @[:@3.2]
  input          clock, // @[:@4.4]
  input          reset, // @[:@5.4]
  input  [162:0] io_a, // @[:@6.4]
  input  [162:0] io_p, // @[:@6.4]
  input          io_bi, // @[:@6.4]
  output [162:0] io_aout, // @[:@6.4]
  output [162:0] io_pout // @[:@6.4]
);
  wire [161:0] _T_15; // @[OneBit.scala 18:24:@8.4]
  wire [162:0] aShift; // @[Cat.scala 30:58:@9.4]
  wire  _T_17; // @[OneBit.scala 19:22:@10.4]
  wire [162:0] _T_27; // @[OneBit.scala 19:44:@14.4]
  wire [162:0] _T_31; // @[OneBit.scala 20:38:@18.4]
  assign _T_15 = io_a[161:0]; // @[OneBit.scala 18:24:@8.4]
  assign aShift = {_T_15,1'h0}; // @[Cat.scala 30:58:@9.4]
  assign _T_17 = io_a[162]; // @[OneBit.scala 19:22:@10.4]
  assign _T_27 = aShift ^ 163'hc9; // @[OneBit.scala 19:44:@14.4]
  assign _T_31 = io_a ^ io_p; // @[OneBit.scala 20:38:@18.4]
  assign io_aout = _T_17 ? _T_27 : aShift; // @[OneBit.scala 19:11:@16.4]
  assign io_pout = io_bi ? _T_31 : io_p; // @[OneBit.scala 20:11:@20.4]
endmodule
