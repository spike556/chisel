module RamSync( // @[:@3.2]
  input          clock, // @[:@4.4]
  input          io_re, // @[:@6.4]
  input          io_we, // @[:@6.4]
  input  [7:0]   io_ra, // @[:@6.4]
  input  [7:0]   io_wa, // @[:@6.4]
  input  [511:0] io_di, // @[:@6.4]
  output [511:0] io_dout // @[:@6.4]
);
  reg [511:0] mem [0:255]; // @[RamSync.scala 26:24:@8.4]
  reg [511:0] _RAND_0;
  wire [511:0] mem__T_23_data; // @[RamSync.scala 26:24:@8.4]
  wire [7:0] mem__T_23_addr; // @[RamSync.scala 26:24:@8.4]
  wire [511:0] mem__T_21_data; // @[RamSync.scala 26:24:@8.4]
  wire [7:0] mem__T_21_addr; // @[RamSync.scala 26:24:@8.4]
  wire  mem__T_21_mask; // @[RamSync.scala 26:24:@8.4]
  wire  mem__T_21_en; // @[RamSync.scala 26:24:@8.4]
  wire [511:0] _GEN_3; // @[RamSync.scala 32:20:@15.6]
  wire  _GEN_12; // @[RamSync.scala 28:16:@9.4]
  reg [7:0] mem__T_23_addr_pipe_0;
  reg [31:0] _RAND_1;
  wire  _GEN_13;
  assign mem__T_23_addr = mem__T_23_addr_pipe_0;
  assign mem__T_23_data = mem[mem__T_23_addr]; // @[RamSync.scala 26:24:@8.4]
  assign mem__T_21_data = io_di;
  assign mem__T_21_addr = io_wa;
  assign mem__T_21_mask = 1'h1;
  assign mem__T_21_en = io_we;
  assign _GEN_3 = io_re ? mem__T_23_data : 512'h0; // @[RamSync.scala 32:20:@15.6]
  assign _GEN_12 = io_we ? 1'h0 : io_re; // @[RamSync.scala 28:16:@9.4]
  assign io_dout = io_we ? 512'h0 : _GEN_3; // @[RamSync.scala 30:13:@12.6 RamSync.scala 33:13:@17.8 RamSync.scala 35:13:@20.8]
  assign _GEN_13 = _GEN_12;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {16{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    mem[initvar] = _RAND_0[511:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem__T_23_addr_pipe_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem__T_21_en & mem__T_21_mask) begin
      mem[mem__T_21_addr] <= mem__T_21_data; // @[RamSync.scala 26:24:@8.4]
    end
    if (_GEN_13) begin
      mem__T_23_addr_pipe_0 <= io_ra;
    end
  end
endmodule
module Cbuf( // @[:@643.2]
  input           clock, // @[:@644.4]
  input           reset, // @[:@645.4]
  input  [31:0]   io_pwrbus_ram_pd, // @[:@646.4]
  input  [1023:0] io_cdma2bufWt_data, // @[:@646.4]
  input  [11:0]   io_cdma2bufWt_addr, // @[:@646.4]
  input           io_cdma2bufWt_enable, // @[:@646.4]
  input  [1:0]    io_cdma2bufWt_hsel, // @[:@646.4]
  input  [1023:0] io_cdma2bufDat_data, // @[:@646.4]
  input  [11:0]   io_cdma2bufDat_addr, // @[:@646.4]
  input           io_cdma2bufDat_enable, // @[:@646.4]
  input  [1:0]    io_cdma2bufDat_hsel, // @[:@646.4]
  input  [11:0]   io_sc2bufDat_addr, // @[:@646.4]
  input           io_sc2bufDat_enable, // @[:@646.4]
  output [1023:0] io_sc2bufDat_data, // @[:@646.4]
  output          io_sc2bufDat_valid, // @[:@646.4]
  input  [11:0]   io_sc2bufWt_addr, // @[:@646.4]
  input           io_sc2bufWt_enable, // @[:@646.4]
  output [1023:0] io_sc2bufWt_data, // @[:@646.4]
  output          io_sc2bufWt_valid, // @[:@646.4]
  input  [11:0]   io_sc2bufWMB_addr, // @[:@646.4]
  input           io_sc2bufWMB_enable, // @[:@646.4]
  output [1023:0] io_sc2bufWMB_data, // @[:@646.4]
  output          io_sc2bufWMB_valid // @[:@646.4]
);
  wire  RamSync_clock; // @[Cbuf.scala 43:52:@648.4]
  wire  RamSync_io_re; // @[Cbuf.scala 43:52:@648.4]
  wire  RamSync_io_we; // @[Cbuf.scala 43:52:@648.4]
  wire [7:0] RamSync_io_ra; // @[Cbuf.scala 43:52:@648.4]
  wire [7:0] RamSync_io_wa; // @[Cbuf.scala 43:52:@648.4]
  wire [511:0] RamSync_io_di; // @[Cbuf.scala 43:52:@648.4]
  wire [511:0] RamSync_io_dout; // @[Cbuf.scala 43:52:@648.4]
  wire  RamSync_1_clock; // @[Cbuf.scala 43:52:@651.4]
  wire  RamSync_1_io_re; // @[Cbuf.scala 43:52:@651.4]
  wire  RamSync_1_io_we; // @[Cbuf.scala 43:52:@651.4]
  wire [7:0] RamSync_1_io_ra; // @[Cbuf.scala 43:52:@651.4]
  wire [7:0] RamSync_1_io_wa; // @[Cbuf.scala 43:52:@651.4]
  wire [511:0] RamSync_1_io_di; // @[Cbuf.scala 43:52:@651.4]
  wire [511:0] RamSync_1_io_dout; // @[Cbuf.scala 43:52:@651.4]
  wire  RamSync_2_clock; // @[Cbuf.scala 43:52:@654.4]
  wire  RamSync_2_io_re; // @[Cbuf.scala 43:52:@654.4]
  wire  RamSync_2_io_we; // @[Cbuf.scala 43:52:@654.4]
  wire [7:0] RamSync_2_io_ra; // @[Cbuf.scala 43:52:@654.4]
  wire [7:0] RamSync_2_io_wa; // @[Cbuf.scala 43:52:@654.4]
  wire [511:0] RamSync_2_io_di; // @[Cbuf.scala 43:52:@654.4]
  wire [511:0] RamSync_2_io_dout; // @[Cbuf.scala 43:52:@654.4]
  wire  RamSync_3_clock; // @[Cbuf.scala 43:52:@657.4]
  wire  RamSync_3_io_re; // @[Cbuf.scala 43:52:@657.4]
  wire  RamSync_3_io_we; // @[Cbuf.scala 43:52:@657.4]
  wire [7:0] RamSync_3_io_ra; // @[Cbuf.scala 43:52:@657.4]
  wire [7:0] RamSync_3_io_wa; // @[Cbuf.scala 43:52:@657.4]
  wire [511:0] RamSync_3_io_di; // @[Cbuf.scala 43:52:@657.4]
  wire [511:0] RamSync_3_io_dout; // @[Cbuf.scala 43:52:@657.4]
  wire  RamSync_4_clock; // @[Cbuf.scala 43:52:@660.4]
  wire  RamSync_4_io_re; // @[Cbuf.scala 43:52:@660.4]
  wire  RamSync_4_io_we; // @[Cbuf.scala 43:52:@660.4]
  wire [7:0] RamSync_4_io_ra; // @[Cbuf.scala 43:52:@660.4]
  wire [7:0] RamSync_4_io_wa; // @[Cbuf.scala 43:52:@660.4]
  wire [511:0] RamSync_4_io_di; // @[Cbuf.scala 43:52:@660.4]
  wire [511:0] RamSync_4_io_dout; // @[Cbuf.scala 43:52:@660.4]
  wire  RamSync_5_clock; // @[Cbuf.scala 43:52:@663.4]
  wire  RamSync_5_io_re; // @[Cbuf.scala 43:52:@663.4]
  wire  RamSync_5_io_we; // @[Cbuf.scala 43:52:@663.4]
  wire [7:0] RamSync_5_io_ra; // @[Cbuf.scala 43:52:@663.4]
  wire [7:0] RamSync_5_io_wa; // @[Cbuf.scala 43:52:@663.4]
  wire [511:0] RamSync_5_io_di; // @[Cbuf.scala 43:52:@663.4]
  wire [511:0] RamSync_5_io_dout; // @[Cbuf.scala 43:52:@663.4]
  wire  RamSync_6_clock; // @[Cbuf.scala 43:52:@666.4]
  wire  RamSync_6_io_re; // @[Cbuf.scala 43:52:@666.4]
  wire  RamSync_6_io_we; // @[Cbuf.scala 43:52:@666.4]
  wire [7:0] RamSync_6_io_ra; // @[Cbuf.scala 43:52:@666.4]
  wire [7:0] RamSync_6_io_wa; // @[Cbuf.scala 43:52:@666.4]
  wire [511:0] RamSync_6_io_di; // @[Cbuf.scala 43:52:@666.4]
  wire [511:0] RamSync_6_io_dout; // @[Cbuf.scala 43:52:@666.4]
  wire  RamSync_7_clock; // @[Cbuf.scala 43:52:@669.4]
  wire  RamSync_7_io_re; // @[Cbuf.scala 43:52:@669.4]
  wire  RamSync_7_io_we; // @[Cbuf.scala 43:52:@669.4]
  wire [7:0] RamSync_7_io_ra; // @[Cbuf.scala 43:52:@669.4]
  wire [7:0] RamSync_7_io_wa; // @[Cbuf.scala 43:52:@669.4]
  wire [511:0] RamSync_7_io_di; // @[Cbuf.scala 43:52:@669.4]
  wire [511:0] RamSync_7_io_dout; // @[Cbuf.scala 43:52:@669.4]
  wire  RamSync_8_clock; // @[Cbuf.scala 43:52:@672.4]
  wire  RamSync_8_io_re; // @[Cbuf.scala 43:52:@672.4]
  wire  RamSync_8_io_we; // @[Cbuf.scala 43:52:@672.4]
  wire [7:0] RamSync_8_io_ra; // @[Cbuf.scala 43:52:@672.4]
  wire [7:0] RamSync_8_io_wa; // @[Cbuf.scala 43:52:@672.4]
  wire [511:0] RamSync_8_io_di; // @[Cbuf.scala 43:52:@672.4]
  wire [511:0] RamSync_8_io_dout; // @[Cbuf.scala 43:52:@672.4]
  wire  RamSync_9_clock; // @[Cbuf.scala 43:52:@675.4]
  wire  RamSync_9_io_re; // @[Cbuf.scala 43:52:@675.4]
  wire  RamSync_9_io_we; // @[Cbuf.scala 43:52:@675.4]
  wire [7:0] RamSync_9_io_ra; // @[Cbuf.scala 43:52:@675.4]
  wire [7:0] RamSync_9_io_wa; // @[Cbuf.scala 43:52:@675.4]
  wire [511:0] RamSync_9_io_di; // @[Cbuf.scala 43:52:@675.4]
  wire [511:0] RamSync_9_io_dout; // @[Cbuf.scala 43:52:@675.4]
  wire  RamSync_10_clock; // @[Cbuf.scala 43:52:@678.4]
  wire  RamSync_10_io_re; // @[Cbuf.scala 43:52:@678.4]
  wire  RamSync_10_io_we; // @[Cbuf.scala 43:52:@678.4]
  wire [7:0] RamSync_10_io_ra; // @[Cbuf.scala 43:52:@678.4]
  wire [7:0] RamSync_10_io_wa; // @[Cbuf.scala 43:52:@678.4]
  wire [511:0] RamSync_10_io_di; // @[Cbuf.scala 43:52:@678.4]
  wire [511:0] RamSync_10_io_dout; // @[Cbuf.scala 43:52:@678.4]
  wire  RamSync_11_clock; // @[Cbuf.scala 43:52:@681.4]
  wire  RamSync_11_io_re; // @[Cbuf.scala 43:52:@681.4]
  wire  RamSync_11_io_we; // @[Cbuf.scala 43:52:@681.4]
  wire [7:0] RamSync_11_io_ra; // @[Cbuf.scala 43:52:@681.4]
  wire [7:0] RamSync_11_io_wa; // @[Cbuf.scala 43:52:@681.4]
  wire [511:0] RamSync_11_io_di; // @[Cbuf.scala 43:52:@681.4]
  wire [511:0] RamSync_11_io_dout; // @[Cbuf.scala 43:52:@681.4]
  wire  RamSync_12_clock; // @[Cbuf.scala 43:52:@684.4]
  wire  RamSync_12_io_re; // @[Cbuf.scala 43:52:@684.4]
  wire  RamSync_12_io_we; // @[Cbuf.scala 43:52:@684.4]
  wire [7:0] RamSync_12_io_ra; // @[Cbuf.scala 43:52:@684.4]
  wire [7:0] RamSync_12_io_wa; // @[Cbuf.scala 43:52:@684.4]
  wire [511:0] RamSync_12_io_di; // @[Cbuf.scala 43:52:@684.4]
  wire [511:0] RamSync_12_io_dout; // @[Cbuf.scala 43:52:@684.4]
  wire  RamSync_13_clock; // @[Cbuf.scala 43:52:@687.4]
  wire  RamSync_13_io_re; // @[Cbuf.scala 43:52:@687.4]
  wire  RamSync_13_io_we; // @[Cbuf.scala 43:52:@687.4]
  wire [7:0] RamSync_13_io_ra; // @[Cbuf.scala 43:52:@687.4]
  wire [7:0] RamSync_13_io_wa; // @[Cbuf.scala 43:52:@687.4]
  wire [511:0] RamSync_13_io_di; // @[Cbuf.scala 43:52:@687.4]
  wire [511:0] RamSync_13_io_dout; // @[Cbuf.scala 43:52:@687.4]
  wire  RamSync_14_clock; // @[Cbuf.scala 43:52:@690.4]
  wire  RamSync_14_io_re; // @[Cbuf.scala 43:52:@690.4]
  wire  RamSync_14_io_we; // @[Cbuf.scala 43:52:@690.4]
  wire [7:0] RamSync_14_io_ra; // @[Cbuf.scala 43:52:@690.4]
  wire [7:0] RamSync_14_io_wa; // @[Cbuf.scala 43:52:@690.4]
  wire [511:0] RamSync_14_io_di; // @[Cbuf.scala 43:52:@690.4]
  wire [511:0] RamSync_14_io_dout; // @[Cbuf.scala 43:52:@690.4]
  wire  RamSync_15_clock; // @[Cbuf.scala 43:52:@693.4]
  wire  RamSync_15_io_re; // @[Cbuf.scala 43:52:@693.4]
  wire  RamSync_15_io_we; // @[Cbuf.scala 43:52:@693.4]
  wire [7:0] RamSync_15_io_ra; // @[Cbuf.scala 43:52:@693.4]
  wire [7:0] RamSync_15_io_wa; // @[Cbuf.scala 43:52:@693.4]
  wire [511:0] RamSync_15_io_di; // @[Cbuf.scala 43:52:@693.4]
  wire [511:0] RamSync_15_io_dout; // @[Cbuf.scala 43:52:@693.4]
  wire  RamSync_16_clock; // @[Cbuf.scala 43:52:@696.4]
  wire  RamSync_16_io_re; // @[Cbuf.scala 43:52:@696.4]
  wire  RamSync_16_io_we; // @[Cbuf.scala 43:52:@696.4]
  wire [7:0] RamSync_16_io_ra; // @[Cbuf.scala 43:52:@696.4]
  wire [7:0] RamSync_16_io_wa; // @[Cbuf.scala 43:52:@696.4]
  wire [511:0] RamSync_16_io_di; // @[Cbuf.scala 43:52:@696.4]
  wire [511:0] RamSync_16_io_dout; // @[Cbuf.scala 43:52:@696.4]
  wire  RamSync_17_clock; // @[Cbuf.scala 43:52:@699.4]
  wire  RamSync_17_io_re; // @[Cbuf.scala 43:52:@699.4]
  wire  RamSync_17_io_we; // @[Cbuf.scala 43:52:@699.4]
  wire [7:0] RamSync_17_io_ra; // @[Cbuf.scala 43:52:@699.4]
  wire [7:0] RamSync_17_io_wa; // @[Cbuf.scala 43:52:@699.4]
  wire [511:0] RamSync_17_io_di; // @[Cbuf.scala 43:52:@699.4]
  wire [511:0] RamSync_17_io_dout; // @[Cbuf.scala 43:52:@699.4]
  wire  RamSync_18_clock; // @[Cbuf.scala 43:52:@702.4]
  wire  RamSync_18_io_re; // @[Cbuf.scala 43:52:@702.4]
  wire  RamSync_18_io_we; // @[Cbuf.scala 43:52:@702.4]
  wire [7:0] RamSync_18_io_ra; // @[Cbuf.scala 43:52:@702.4]
  wire [7:0] RamSync_18_io_wa; // @[Cbuf.scala 43:52:@702.4]
  wire [511:0] RamSync_18_io_di; // @[Cbuf.scala 43:52:@702.4]
  wire [511:0] RamSync_18_io_dout; // @[Cbuf.scala 43:52:@702.4]
  wire  RamSync_19_clock; // @[Cbuf.scala 43:52:@705.4]
  wire  RamSync_19_io_re; // @[Cbuf.scala 43:52:@705.4]
  wire  RamSync_19_io_we; // @[Cbuf.scala 43:52:@705.4]
  wire [7:0] RamSync_19_io_ra; // @[Cbuf.scala 43:52:@705.4]
  wire [7:0] RamSync_19_io_wa; // @[Cbuf.scala 43:52:@705.4]
  wire [511:0] RamSync_19_io_di; // @[Cbuf.scala 43:52:@705.4]
  wire [511:0] RamSync_19_io_dout; // @[Cbuf.scala 43:52:@705.4]
  wire  RamSync_20_clock; // @[Cbuf.scala 43:52:@708.4]
  wire  RamSync_20_io_re; // @[Cbuf.scala 43:52:@708.4]
  wire  RamSync_20_io_we; // @[Cbuf.scala 43:52:@708.4]
  wire [7:0] RamSync_20_io_ra; // @[Cbuf.scala 43:52:@708.4]
  wire [7:0] RamSync_20_io_wa; // @[Cbuf.scala 43:52:@708.4]
  wire [511:0] RamSync_20_io_di; // @[Cbuf.scala 43:52:@708.4]
  wire [511:0] RamSync_20_io_dout; // @[Cbuf.scala 43:52:@708.4]
  wire  RamSync_21_clock; // @[Cbuf.scala 43:52:@711.4]
  wire  RamSync_21_io_re; // @[Cbuf.scala 43:52:@711.4]
  wire  RamSync_21_io_we; // @[Cbuf.scala 43:52:@711.4]
  wire [7:0] RamSync_21_io_ra; // @[Cbuf.scala 43:52:@711.4]
  wire [7:0] RamSync_21_io_wa; // @[Cbuf.scala 43:52:@711.4]
  wire [511:0] RamSync_21_io_di; // @[Cbuf.scala 43:52:@711.4]
  wire [511:0] RamSync_21_io_dout; // @[Cbuf.scala 43:52:@711.4]
  wire  RamSync_22_clock; // @[Cbuf.scala 43:52:@714.4]
  wire  RamSync_22_io_re; // @[Cbuf.scala 43:52:@714.4]
  wire  RamSync_22_io_we; // @[Cbuf.scala 43:52:@714.4]
  wire [7:0] RamSync_22_io_ra; // @[Cbuf.scala 43:52:@714.4]
  wire [7:0] RamSync_22_io_wa; // @[Cbuf.scala 43:52:@714.4]
  wire [511:0] RamSync_22_io_di; // @[Cbuf.scala 43:52:@714.4]
  wire [511:0] RamSync_22_io_dout; // @[Cbuf.scala 43:52:@714.4]
  wire  RamSync_23_clock; // @[Cbuf.scala 43:52:@717.4]
  wire  RamSync_23_io_re; // @[Cbuf.scala 43:52:@717.4]
  wire  RamSync_23_io_we; // @[Cbuf.scala 43:52:@717.4]
  wire [7:0] RamSync_23_io_ra; // @[Cbuf.scala 43:52:@717.4]
  wire [7:0] RamSync_23_io_wa; // @[Cbuf.scala 43:52:@717.4]
  wire [511:0] RamSync_23_io_di; // @[Cbuf.scala 43:52:@717.4]
  wire [511:0] RamSync_23_io_dout; // @[Cbuf.scala 43:52:@717.4]
  wire  RamSync_24_clock; // @[Cbuf.scala 43:52:@720.4]
  wire  RamSync_24_io_re; // @[Cbuf.scala 43:52:@720.4]
  wire  RamSync_24_io_we; // @[Cbuf.scala 43:52:@720.4]
  wire [7:0] RamSync_24_io_ra; // @[Cbuf.scala 43:52:@720.4]
  wire [7:0] RamSync_24_io_wa; // @[Cbuf.scala 43:52:@720.4]
  wire [511:0] RamSync_24_io_di; // @[Cbuf.scala 43:52:@720.4]
  wire [511:0] RamSync_24_io_dout; // @[Cbuf.scala 43:52:@720.4]
  wire  RamSync_25_clock; // @[Cbuf.scala 43:52:@723.4]
  wire  RamSync_25_io_re; // @[Cbuf.scala 43:52:@723.4]
  wire  RamSync_25_io_we; // @[Cbuf.scala 43:52:@723.4]
  wire [7:0] RamSync_25_io_ra; // @[Cbuf.scala 43:52:@723.4]
  wire [7:0] RamSync_25_io_wa; // @[Cbuf.scala 43:52:@723.4]
  wire [511:0] RamSync_25_io_di; // @[Cbuf.scala 43:52:@723.4]
  wire [511:0] RamSync_25_io_dout; // @[Cbuf.scala 43:52:@723.4]
  wire  RamSync_26_clock; // @[Cbuf.scala 43:52:@726.4]
  wire  RamSync_26_io_re; // @[Cbuf.scala 43:52:@726.4]
  wire  RamSync_26_io_we; // @[Cbuf.scala 43:52:@726.4]
  wire [7:0] RamSync_26_io_ra; // @[Cbuf.scala 43:52:@726.4]
  wire [7:0] RamSync_26_io_wa; // @[Cbuf.scala 43:52:@726.4]
  wire [511:0] RamSync_26_io_di; // @[Cbuf.scala 43:52:@726.4]
  wire [511:0] RamSync_26_io_dout; // @[Cbuf.scala 43:52:@726.4]
  wire  RamSync_27_clock; // @[Cbuf.scala 43:52:@729.4]
  wire  RamSync_27_io_re; // @[Cbuf.scala 43:52:@729.4]
  wire  RamSync_27_io_we; // @[Cbuf.scala 43:52:@729.4]
  wire [7:0] RamSync_27_io_ra; // @[Cbuf.scala 43:52:@729.4]
  wire [7:0] RamSync_27_io_wa; // @[Cbuf.scala 43:52:@729.4]
  wire [511:0] RamSync_27_io_di; // @[Cbuf.scala 43:52:@729.4]
  wire [511:0] RamSync_27_io_dout; // @[Cbuf.scala 43:52:@729.4]
  wire  RamSync_28_clock; // @[Cbuf.scala 43:52:@732.4]
  wire  RamSync_28_io_re; // @[Cbuf.scala 43:52:@732.4]
  wire  RamSync_28_io_we; // @[Cbuf.scala 43:52:@732.4]
  wire [7:0] RamSync_28_io_ra; // @[Cbuf.scala 43:52:@732.4]
  wire [7:0] RamSync_28_io_wa; // @[Cbuf.scala 43:52:@732.4]
  wire [511:0] RamSync_28_io_di; // @[Cbuf.scala 43:52:@732.4]
  wire [511:0] RamSync_28_io_dout; // @[Cbuf.scala 43:52:@732.4]
  wire  RamSync_29_clock; // @[Cbuf.scala 43:52:@735.4]
  wire  RamSync_29_io_re; // @[Cbuf.scala 43:52:@735.4]
  wire  RamSync_29_io_we; // @[Cbuf.scala 43:52:@735.4]
  wire [7:0] RamSync_29_io_ra; // @[Cbuf.scala 43:52:@735.4]
  wire [7:0] RamSync_29_io_wa; // @[Cbuf.scala 43:52:@735.4]
  wire [511:0] RamSync_29_io_di; // @[Cbuf.scala 43:52:@735.4]
  wire [511:0] RamSync_29_io_dout; // @[Cbuf.scala 43:52:@735.4]
  wire  RamSync_30_clock; // @[Cbuf.scala 43:52:@738.4]
  wire  RamSync_30_io_re; // @[Cbuf.scala 43:52:@738.4]
  wire  RamSync_30_io_we; // @[Cbuf.scala 43:52:@738.4]
  wire [7:0] RamSync_30_io_ra; // @[Cbuf.scala 43:52:@738.4]
  wire [7:0] RamSync_30_io_wa; // @[Cbuf.scala 43:52:@738.4]
  wire [511:0] RamSync_30_io_di; // @[Cbuf.scala 43:52:@738.4]
  wire [511:0] RamSync_30_io_dout; // @[Cbuf.scala 43:52:@738.4]
  wire  RamSync_31_clock; // @[Cbuf.scala 43:52:@741.4]
  wire  RamSync_31_io_re; // @[Cbuf.scala 43:52:@741.4]
  wire  RamSync_31_io_we; // @[Cbuf.scala 43:52:@741.4]
  wire [7:0] RamSync_31_io_ra; // @[Cbuf.scala 43:52:@741.4]
  wire [7:0] RamSync_31_io_wa; // @[Cbuf.scala 43:52:@741.4]
  wire [511:0] RamSync_31_io_di; // @[Cbuf.scala 43:52:@741.4]
  wire [511:0] RamSync_31_io_dout; // @[Cbuf.scala 43:52:@741.4]
  wire [3:0] _T_1533; // @[Cbuf.scala 54:30:@906.4]
  wire  _T_1558; // @[Cbuf.scala 54:87:@907.4]
  wire  _T_1559; // @[Cbuf.scala 54:66:@908.4]
  wire  datWreq_0_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_1_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_2_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_3_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_4_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_5_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_6_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_7_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_8_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_9_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_10_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_11_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_12_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_13_0; // @[Cbuf.scala 54:41:@909.4]
  wire  datWreq_14_0; // @[Cbuf.scala 54:41:@909.4]
  wire  _T_1585; // @[Cbuf.scala 55:87:@911.4]
  wire  _T_1586; // @[Cbuf.scala 55:66:@912.4]
  wire  datWreq_0_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_1_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_2_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_3_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_4_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_5_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_6_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_7_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_8_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_9_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_10_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_11_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_12_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_13_1; // @[Cbuf.scala 55:41:@913.4]
  wire  datWreq_14_1; // @[Cbuf.scala 55:41:@913.4]
  wire [3:0] _T_1587; // @[Cbuf.scala 58:28:@914.4]
  wire  _T_1612; // @[Cbuf.scala 58:85:@915.4]
  wire  _T_1614; // @[Cbuf.scala 58:66:@916.4]
  wire  _T_1615; // @[Cbuf.scala 58:63:@917.4]
  wire  wtWreq_1_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_2_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_3_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_4_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_5_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_6_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_7_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_8_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_9_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_10_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_11_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_12_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_13_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_14_0; // @[Cbuf.scala 58:39:@918.4]
  wire  wtWreq_15_0; // @[Cbuf.scala 58:39:@918.4]
  wire  _T_1642; // @[Cbuf.scala 59:63:@921.4]
  wire  wtWreq_1_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_2_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_3_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_4_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_5_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_6_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_7_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_8_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_9_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_10_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_11_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_12_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_13_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_14_1; // @[Cbuf.scala 59:39:@922.4]
  wire  wtWreq_15_1; // @[Cbuf.scala 59:39:@922.4]
  reg  ramWreqd1_0_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_0;
  reg  ramWreqd1_0_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_1;
  reg  ramWreqd1_1_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_2;
  reg  ramWreqd1_1_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_3;
  reg  ramWreqd1_2_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_4;
  reg  ramWreqd1_2_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_5;
  reg  ramWreqd1_3_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_6;
  reg  ramWreqd1_3_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_7;
  reg  ramWreqd1_4_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_8;
  reg  ramWreqd1_4_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_9;
  reg  ramWreqd1_5_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_10;
  reg  ramWreqd1_5_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_11;
  reg  ramWreqd1_6_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_12;
  reg  ramWreqd1_6_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_13;
  reg  ramWreqd1_7_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_14;
  reg  ramWreqd1_7_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_15;
  reg  ramWreqd1_8_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_16;
  reg  ramWreqd1_8_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_17;
  reg  ramWreqd1_9_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_18;
  reg  ramWreqd1_9_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_19;
  reg  ramWreqd1_10_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_20;
  reg  ramWreqd1_10_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_21;
  reg  ramWreqd1_11_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_22;
  reg  ramWreqd1_11_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_23;
  reg  ramWreqd1_12_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_24;
  reg  ramWreqd1_12_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_25;
  reg  ramWreqd1_13_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_26;
  reg  ramWreqd1_13_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_27;
  reg  ramWreqd1_14_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_28;
  reg  ramWreqd1_14_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_29;
  reg  ramWreqd1_15_0; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_30;
  reg  ramWreqd1_15_1; // @[Cbuf.scala 64:26:@1004.4]
  reg [31:0] _RAND_31;
  reg [7:0] ramp0Addrd1; // @[Cbuf.scala 65:28:@1006.4]
  reg [31:0] _RAND_32;
  reg [7:0] ramp1Addrd1; // @[Cbuf.scala 66:28:@1009.4]
  reg [31:0] _RAND_33;
  reg [511:0] ramp0DatLod1; // @[Cbuf.scala 67:29:@1012.4]
  reg [511:0] _RAND_34;
  reg [511:0] ramp0DatHid1; // @[Cbuf.scala 68:29:@1015.4]
  reg [511:0] _RAND_35;
  reg [511:0] ramp1WtLod1; // @[Cbuf.scala 69:28:@1018.4]
  reg [511:0] _RAND_36;
  reg [511:0] ramp1WtHid1; // @[Cbuf.scala 70:28:@1021.4]
  reg [511:0] _RAND_37;
  wire  _T_4142; // @[Cbuf.scala 84:40:@1025.4]
  wire  _T_4143; // @[Cbuf.scala 85:40:@1027.4]
  wire  _T_4144; // @[Cbuf.scala 84:40:@1029.4]
  wire  _T_4145; // @[Cbuf.scala 85:40:@1031.4]
  wire  _T_4146; // @[Cbuf.scala 84:40:@1033.4]
  wire  _T_4147; // @[Cbuf.scala 85:40:@1035.4]
  wire  _T_4148; // @[Cbuf.scala 84:40:@1037.4]
  wire  _T_4149; // @[Cbuf.scala 85:40:@1039.4]
  wire  _T_4150; // @[Cbuf.scala 84:40:@1041.4]
  wire  _T_4151; // @[Cbuf.scala 85:40:@1043.4]
  wire  _T_4152; // @[Cbuf.scala 84:40:@1045.4]
  wire  _T_4153; // @[Cbuf.scala 85:40:@1047.4]
  wire  _T_4154; // @[Cbuf.scala 84:40:@1049.4]
  wire  _T_4155; // @[Cbuf.scala 85:40:@1051.4]
  wire  _T_4156; // @[Cbuf.scala 84:40:@1053.4]
  wire  _T_4157; // @[Cbuf.scala 85:40:@1055.4]
  wire  _T_4158; // @[Cbuf.scala 84:40:@1057.4]
  wire  _T_4159; // @[Cbuf.scala 85:40:@1059.4]
  wire  _T_4160; // @[Cbuf.scala 84:40:@1061.4]
  wire  _T_4161; // @[Cbuf.scala 85:40:@1063.4]
  wire  _T_4162; // @[Cbuf.scala 84:40:@1065.4]
  wire  _T_4163; // @[Cbuf.scala 85:40:@1067.4]
  wire  _T_4164; // @[Cbuf.scala 84:40:@1069.4]
  wire  _T_4165; // @[Cbuf.scala 85:40:@1071.4]
  wire  _T_4166; // @[Cbuf.scala 84:40:@1073.4]
  wire  _T_4167; // @[Cbuf.scala 85:40:@1075.4]
  wire  _T_4168; // @[Cbuf.scala 84:40:@1077.4]
  wire  _T_4169; // @[Cbuf.scala 85:40:@1079.4]
  wire [7:0] _T_5162; // @[Cbuf.scala 105:31:@1465.4]
  wire [7:0] _T_5166; // @[Cbuf.scala 105:80:@1467.4]
  wire [7:0] _T_5171; // @[Cbuf.scala 106:31:@1471.4]
  wire [7:0] _T_5175; // @[Cbuf.scala 106:80:@1473.4]
  wire [511:0] _T_5180; // @[Cbuf.scala 107:31:@1477.4]
  wire [511:0] _T_5184; // @[Cbuf.scala 107:81:@1479.4]
  wire [511:0] _T_5189; // @[Cbuf.scala 108:31:@1483.4]
  wire [511:0] _T_5193; // @[Cbuf.scala 108:81:@1485.4]
  wire [7:0] _T_5198; // @[Cbuf.scala 105:31:@1489.4]
  wire [7:0] _T_5202; // @[Cbuf.scala 105:80:@1491.4]
  wire [7:0] _T_5207; // @[Cbuf.scala 106:31:@1495.4]
  wire [7:0] _T_5211; // @[Cbuf.scala 106:80:@1497.4]
  wire [511:0] _T_5216; // @[Cbuf.scala 107:31:@1501.4]
  wire [511:0] _T_5220; // @[Cbuf.scala 107:81:@1503.4]
  wire [511:0] _T_5225; // @[Cbuf.scala 108:31:@1507.4]
  wire [511:0] _T_5229; // @[Cbuf.scala 108:81:@1509.4]
  wire [7:0] _T_5234; // @[Cbuf.scala 105:31:@1513.4]
  wire [7:0] _T_5238; // @[Cbuf.scala 105:80:@1515.4]
  wire [7:0] _T_5243; // @[Cbuf.scala 106:31:@1519.4]
  wire [7:0] _T_5247; // @[Cbuf.scala 106:80:@1521.4]
  wire [511:0] _T_5252; // @[Cbuf.scala 107:31:@1525.4]
  wire [511:0] _T_5256; // @[Cbuf.scala 107:81:@1527.4]
  wire [511:0] _T_5261; // @[Cbuf.scala 108:31:@1531.4]
  wire [511:0] _T_5265; // @[Cbuf.scala 108:81:@1533.4]
  wire [7:0] _T_5270; // @[Cbuf.scala 105:31:@1537.4]
  wire [7:0] _T_5274; // @[Cbuf.scala 105:80:@1539.4]
  wire [7:0] _T_5279; // @[Cbuf.scala 106:31:@1543.4]
  wire [7:0] _T_5283; // @[Cbuf.scala 106:80:@1545.4]
  wire [511:0] _T_5288; // @[Cbuf.scala 107:31:@1549.4]
  wire [511:0] _T_5292; // @[Cbuf.scala 107:81:@1551.4]
  wire [511:0] _T_5297; // @[Cbuf.scala 108:31:@1555.4]
  wire [511:0] _T_5301; // @[Cbuf.scala 108:81:@1557.4]
  wire [7:0] _T_5306; // @[Cbuf.scala 105:31:@1561.4]
  wire [7:0] _T_5310; // @[Cbuf.scala 105:80:@1563.4]
  wire [7:0] _T_5315; // @[Cbuf.scala 106:31:@1567.4]
  wire [7:0] _T_5319; // @[Cbuf.scala 106:80:@1569.4]
  wire [511:0] _T_5324; // @[Cbuf.scala 107:31:@1573.4]
  wire [511:0] _T_5328; // @[Cbuf.scala 107:81:@1575.4]
  wire [511:0] _T_5333; // @[Cbuf.scala 108:31:@1579.4]
  wire [511:0] _T_5337; // @[Cbuf.scala 108:81:@1581.4]
  wire [7:0] _T_5342; // @[Cbuf.scala 105:31:@1585.4]
  wire [7:0] _T_5346; // @[Cbuf.scala 105:80:@1587.4]
  wire [7:0] _T_5351; // @[Cbuf.scala 106:31:@1591.4]
  wire [7:0] _T_5355; // @[Cbuf.scala 106:80:@1593.4]
  wire [511:0] _T_5360; // @[Cbuf.scala 107:31:@1597.4]
  wire [511:0] _T_5364; // @[Cbuf.scala 107:81:@1599.4]
  wire [511:0] _T_5369; // @[Cbuf.scala 108:31:@1603.4]
  wire [511:0] _T_5373; // @[Cbuf.scala 108:81:@1605.4]
  wire [7:0] _T_5378; // @[Cbuf.scala 105:31:@1609.4]
  wire [7:0] _T_5382; // @[Cbuf.scala 105:80:@1611.4]
  wire [7:0] _T_5387; // @[Cbuf.scala 106:31:@1615.4]
  wire [7:0] _T_5391; // @[Cbuf.scala 106:80:@1617.4]
  wire [511:0] _T_5396; // @[Cbuf.scala 107:31:@1621.4]
  wire [511:0] _T_5400; // @[Cbuf.scala 107:81:@1623.4]
  wire [511:0] _T_5405; // @[Cbuf.scala 108:31:@1627.4]
  wire [511:0] _T_5409; // @[Cbuf.scala 108:81:@1629.4]
  wire [7:0] _T_5414; // @[Cbuf.scala 105:31:@1633.4]
  wire [7:0] _T_5418; // @[Cbuf.scala 105:80:@1635.4]
  wire [7:0] _T_5423; // @[Cbuf.scala 106:31:@1639.4]
  wire [7:0] _T_5427; // @[Cbuf.scala 106:80:@1641.4]
  wire [511:0] _T_5432; // @[Cbuf.scala 107:31:@1645.4]
  wire [511:0] _T_5436; // @[Cbuf.scala 107:81:@1647.4]
  wire [511:0] _T_5441; // @[Cbuf.scala 108:31:@1651.4]
  wire [511:0] _T_5445; // @[Cbuf.scala 108:81:@1653.4]
  wire [7:0] _T_5450; // @[Cbuf.scala 105:31:@1657.4]
  wire [7:0] _T_5454; // @[Cbuf.scala 105:80:@1659.4]
  wire [7:0] _T_5459; // @[Cbuf.scala 106:31:@1663.4]
  wire [7:0] _T_5463; // @[Cbuf.scala 106:80:@1665.4]
  wire [511:0] _T_5468; // @[Cbuf.scala 107:31:@1669.4]
  wire [511:0] _T_5472; // @[Cbuf.scala 107:81:@1671.4]
  wire [511:0] _T_5477; // @[Cbuf.scala 108:31:@1675.4]
  wire [511:0] _T_5481; // @[Cbuf.scala 108:81:@1677.4]
  wire [7:0] _T_5486; // @[Cbuf.scala 105:31:@1681.4]
  wire [7:0] _T_5490; // @[Cbuf.scala 105:80:@1683.4]
  wire [7:0] _T_5495; // @[Cbuf.scala 106:31:@1687.4]
  wire [7:0] _T_5499; // @[Cbuf.scala 106:80:@1689.4]
  wire [511:0] _T_5504; // @[Cbuf.scala 107:31:@1693.4]
  wire [511:0] _T_5508; // @[Cbuf.scala 107:81:@1695.4]
  wire [511:0] _T_5513; // @[Cbuf.scala 108:31:@1699.4]
  wire [511:0] _T_5517; // @[Cbuf.scala 108:81:@1701.4]
  wire [7:0] _T_5522; // @[Cbuf.scala 105:31:@1705.4]
  wire [7:0] _T_5526; // @[Cbuf.scala 105:80:@1707.4]
  wire [7:0] _T_5531; // @[Cbuf.scala 106:31:@1711.4]
  wire [7:0] _T_5535; // @[Cbuf.scala 106:80:@1713.4]
  wire [511:0] _T_5540; // @[Cbuf.scala 107:31:@1717.4]
  wire [511:0] _T_5544; // @[Cbuf.scala 107:81:@1719.4]
  wire [511:0] _T_5549; // @[Cbuf.scala 108:31:@1723.4]
  wire [511:0] _T_5553; // @[Cbuf.scala 108:81:@1725.4]
  wire [7:0] _T_5558; // @[Cbuf.scala 105:31:@1729.4]
  wire [7:0] _T_5562; // @[Cbuf.scala 105:80:@1731.4]
  wire [7:0] _T_5567; // @[Cbuf.scala 106:31:@1735.4]
  wire [7:0] _T_5571; // @[Cbuf.scala 106:80:@1737.4]
  wire [511:0] _T_5576; // @[Cbuf.scala 107:31:@1741.4]
  wire [511:0] _T_5580; // @[Cbuf.scala 107:81:@1743.4]
  wire [511:0] _T_5585; // @[Cbuf.scala 108:31:@1747.4]
  wire [511:0] _T_5589; // @[Cbuf.scala 108:81:@1749.4]
  wire [7:0] _T_5594; // @[Cbuf.scala 105:31:@1753.4]
  wire [7:0] _T_5598; // @[Cbuf.scala 105:80:@1755.4]
  wire [7:0] _T_5603; // @[Cbuf.scala 106:31:@1759.4]
  wire [7:0] _T_5607; // @[Cbuf.scala 106:80:@1761.4]
  wire [511:0] _T_5612; // @[Cbuf.scala 107:31:@1765.4]
  wire [511:0] _T_5616; // @[Cbuf.scala 107:81:@1767.4]
  wire [511:0] _T_5621; // @[Cbuf.scala 108:31:@1771.4]
  wire [511:0] _T_5625; // @[Cbuf.scala 108:81:@1773.4]
  wire [7:0] _T_5630; // @[Cbuf.scala 105:31:@1777.4]
  wire [7:0] _T_5634; // @[Cbuf.scala 105:80:@1779.4]
  wire [7:0] _T_5639; // @[Cbuf.scala 106:31:@1783.4]
  wire [7:0] _T_5643; // @[Cbuf.scala 106:80:@1785.4]
  wire [511:0] _T_5648; // @[Cbuf.scala 107:31:@1789.4]
  wire [511:0] _T_5652; // @[Cbuf.scala 107:81:@1791.4]
  wire [511:0] _T_5657; // @[Cbuf.scala 108:31:@1795.4]
  wire [511:0] _T_5661; // @[Cbuf.scala 108:81:@1797.4]
  reg  ramWreqd2_0_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_38;
  reg  ramWreqd2_0_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_39;
  reg  ramWreqd2_1_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_40;
  reg  ramWreqd2_1_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_41;
  reg  ramWreqd2_2_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_42;
  reg  ramWreqd2_2_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_43;
  reg  ramWreqd2_3_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_44;
  reg  ramWreqd2_3_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_45;
  reg  ramWreqd2_4_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_46;
  reg  ramWreqd2_4_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_47;
  reg  ramWreqd2_5_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_48;
  reg  ramWreqd2_5_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_49;
  reg  ramWreqd2_6_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_50;
  reg  ramWreqd2_6_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_51;
  reg  ramWreqd2_7_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_52;
  reg  ramWreqd2_7_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_53;
  reg  ramWreqd2_8_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_54;
  reg  ramWreqd2_8_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_55;
  reg  ramWreqd2_9_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_56;
  reg  ramWreqd2_9_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_57;
  reg  ramWreqd2_10_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_58;
  reg  ramWreqd2_10_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_59;
  reg  ramWreqd2_11_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_60;
  reg  ramWreqd2_11_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_61;
  reg  ramWreqd2_12_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_62;
  reg  ramWreqd2_12_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_63;
  reg  ramWreqd2_13_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_64;
  reg  ramWreqd2_13_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_65;
  reg  ramWreqd2_14_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_66;
  reg  ramWreqd2_14_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_67;
  reg  ramWreqd2_15_0; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_68;
  reg  ramWreqd2_15_1; // @[Cbuf.scala 113:26:@1893.4]
  reg [31:0] _RAND_69;
  wire [3:0] _T_10644; // @[Cbuf.scala 129:28:@2524.4]
  wire  datRreq_0_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_1_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_2_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_3_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_4_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_5_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_6_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_7_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_8_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_9_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_10_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_11_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_12_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_13_0; // @[Cbuf.scala 129:36:@2528.4]
  wire  datRreq_14_0; // @[Cbuf.scala 129:36:@2528.4]
  wire [3:0] _T_10687; // @[Cbuf.scala 132:26:@2535.4]
  wire  wtRreq_1_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_2_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_3_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_4_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_5_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_6_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_7_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_8_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_9_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_10_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_11_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_12_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_13_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_14_0; // @[Cbuf.scala 132:34:@2539.4]
  wire  wtRreq_15_0; // @[Cbuf.scala 132:34:@2539.4]
  reg  ramRreq_0_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_70;
  reg  ramRreq_0_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_71;
  reg  ramRreq_1_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_72;
  reg  ramRreq_1_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_73;
  reg  ramRreq_2_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_74;
  reg  ramRreq_2_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_75;
  reg  ramRreq_3_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_76;
  reg  ramRreq_3_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_77;
  reg  ramRreq_4_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_78;
  reg  ramRreq_4_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_79;
  reg  ramRreq_5_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_80;
  reg  ramRreq_5_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_81;
  reg  ramRreq_6_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_82;
  reg  ramRreq_6_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_83;
  reg  ramRreq_7_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_84;
  reg  ramRreq_7_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_85;
  reg  ramRreq_8_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_86;
  reg  ramRreq_8_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_87;
  reg  ramRreq_9_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_88;
  reg  ramRreq_9_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_89;
  reg  ramRreq_10_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_90;
  reg  ramRreq_10_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_91;
  reg  ramRreq_11_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_92;
  reg  ramRreq_11_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_93;
  reg  ramRreq_12_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_94;
  reg  ramRreq_12_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_95;
  reg  ramRreq_13_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_96;
  reg  ramRreq_13_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_97;
  reg  ramRreq_14_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_98;
  reg  ramRreq_14_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_99;
  reg  ramRreq_15_0; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_100;
  reg  ramRreq_15_1; // @[Cbuf.scala 137:24:@2627.4]
  reg [31:0] _RAND_101;
  reg [7:0] ramRaddr_0_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_102;
  reg [7:0] ramRaddr_0_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_103;
  reg [7:0] ramRaddr_1_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_104;
  reg [7:0] ramRaddr_1_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_105;
  reg [7:0] ramRaddr_2_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_106;
  reg [7:0] ramRaddr_2_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_107;
  reg [7:0] ramRaddr_3_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_108;
  reg [7:0] ramRaddr_3_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_109;
  reg [7:0] ramRaddr_4_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_110;
  reg [7:0] ramRaddr_4_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_111;
  reg [7:0] ramRaddr_5_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_112;
  reg [7:0] ramRaddr_5_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_113;
  reg [7:0] ramRaddr_6_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_114;
  reg [7:0] ramRaddr_6_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_115;
  reg [7:0] ramRaddr_7_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_116;
  reg [7:0] ramRaddr_7_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_117;
  reg [7:0] ramRaddr_8_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_118;
  reg [7:0] ramRaddr_8_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_119;
  reg [7:0] ramRaddr_9_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_120;
  reg [7:0] ramRaddr_9_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_121;
  reg [7:0] ramRaddr_10_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_122;
  reg [7:0] ramRaddr_10_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_123;
  reg [7:0] ramRaddr_11_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_124;
  reg [7:0] ramRaddr_11_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_125;
  reg [7:0] ramRaddr_12_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_126;
  reg [7:0] ramRaddr_12_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_127;
  reg [7:0] ramRaddr_13_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_128;
  reg [7:0] ramRaddr_13_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_129;
  reg [7:0] ramRaddr_14_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_130;
  reg [7:0] ramRaddr_14_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_131;
  reg [7:0] ramRaddr_15_0; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_132;
  reg [7:0] ramRaddr_15_1; // @[Cbuf.scala 138:25:@2709.4]
  reg [31:0] _RAND_133;
  wire  _T_15704; // @[Cbuf.scala 149:38:@2712.4]
  wire  _T_15706; // @[Cbuf.scala 149:38:@2716.4]
  wire  _T_15708; // @[Cbuf.scala 149:38:@2720.4]
  wire  _T_15710; // @[Cbuf.scala 149:38:@2724.4]
  wire  _T_15712; // @[Cbuf.scala 149:38:@2728.4]
  wire  _T_15714; // @[Cbuf.scala 149:38:@2732.4]
  wire  _T_15716; // @[Cbuf.scala 149:38:@2736.4]
  wire  _T_15718; // @[Cbuf.scala 149:38:@2740.4]
  wire  _T_15720; // @[Cbuf.scala 149:38:@2744.4]
  wire  _T_15722; // @[Cbuf.scala 149:38:@2748.4]
  wire  _T_15724; // @[Cbuf.scala 149:38:@2752.4]
  wire  _T_15726; // @[Cbuf.scala 149:38:@2756.4]
  wire  _T_15728; // @[Cbuf.scala 149:38:@2760.4]
  wire  _T_15730; // @[Cbuf.scala 149:38:@2764.4]
  wire  _T_15732; // @[Cbuf.scala 145:37:@2768.4]
  wire [11:0] _T_15737; // @[Cbuf.scala 156:28:@2773.4]
  wire [11:0] _T_15745; // @[Cbuf.scala 164:28:@2779.4]
  wire [11:0] _T_15749; // @[Cbuf.scala 164:81:@2781.4]
  wire [11:0] _T_15750; // @[Cbuf.scala 164:76:@2782.4]
  wire [11:0] _T_15763; // @[Cbuf.scala 164:28:@2791.4]
  wire [11:0] _T_15767; // @[Cbuf.scala 164:81:@2793.4]
  wire [11:0] _T_15768; // @[Cbuf.scala 164:76:@2794.4]
  wire [11:0] _T_15781; // @[Cbuf.scala 164:28:@2803.4]
  wire [11:0] _T_15785; // @[Cbuf.scala 164:81:@2805.4]
  wire [11:0] _T_15786; // @[Cbuf.scala 164:76:@2806.4]
  wire [11:0] _T_15799; // @[Cbuf.scala 164:28:@2815.4]
  wire [11:0] _T_15803; // @[Cbuf.scala 164:81:@2817.4]
  wire [11:0] _T_15804; // @[Cbuf.scala 164:76:@2818.4]
  wire [11:0] _T_15817; // @[Cbuf.scala 164:28:@2827.4]
  wire [11:0] _T_15821; // @[Cbuf.scala 164:81:@2829.4]
  wire [11:0] _T_15822; // @[Cbuf.scala 164:76:@2830.4]
  wire [11:0] _T_15835; // @[Cbuf.scala 164:28:@2839.4]
  wire [11:0] _T_15839; // @[Cbuf.scala 164:81:@2841.4]
  wire [11:0] _T_15840; // @[Cbuf.scala 164:76:@2842.4]
  wire [11:0] _T_15853; // @[Cbuf.scala 164:28:@2851.4]
  wire [11:0] _T_15857; // @[Cbuf.scala 164:81:@2853.4]
  wire [11:0] _T_15858; // @[Cbuf.scala 164:76:@2854.4]
  wire [11:0] _T_15871; // @[Cbuf.scala 164:28:@2863.4]
  wire [11:0] _T_15875; // @[Cbuf.scala 164:81:@2865.4]
  wire [11:0] _T_15876; // @[Cbuf.scala 164:76:@2866.4]
  wire [11:0] _T_15889; // @[Cbuf.scala 164:28:@2875.4]
  wire [11:0] _T_15893; // @[Cbuf.scala 164:81:@2877.4]
  wire [11:0] _T_15894; // @[Cbuf.scala 164:76:@2878.4]
  wire [11:0] _T_15907; // @[Cbuf.scala 164:28:@2887.4]
  wire [11:0] _T_15911; // @[Cbuf.scala 164:81:@2889.4]
  wire [11:0] _T_15912; // @[Cbuf.scala 164:76:@2890.4]
  wire [11:0] _T_15925; // @[Cbuf.scala 164:28:@2899.4]
  wire [11:0] _T_15929; // @[Cbuf.scala 164:81:@2901.4]
  wire [11:0] _T_15930; // @[Cbuf.scala 164:76:@2902.4]
  wire [11:0] _T_15943; // @[Cbuf.scala 164:28:@2911.4]
  wire [11:0] _T_15947; // @[Cbuf.scala 164:81:@2913.4]
  wire [11:0] _T_15948; // @[Cbuf.scala 164:76:@2914.4]
  wire [11:0] _T_15961; // @[Cbuf.scala 164:28:@2923.4]
  wire [11:0] _T_15965; // @[Cbuf.scala 164:81:@2925.4]
  wire [11:0] _T_15966; // @[Cbuf.scala 164:76:@2926.4]
  wire [11:0] _T_15979; // @[Cbuf.scala 164:28:@2935.4]
  wire [11:0] _T_15983; // @[Cbuf.scala 164:81:@2937.4]
  wire [11:0] _T_15984; // @[Cbuf.scala 164:76:@2938.4]
  wire [11:0] _T_15997; // @[Cbuf.scala 160:28:@2947.4]
  wire [11:0] _T_16001; // @[Cbuf.scala 160:79:@2949.4]
  wire [11:0] _T_16002; // @[Cbuf.scala 160:74:@2950.4]
  reg  _T_16712_0_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_134;
  reg  _T_16712_0_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_135;
  reg  _T_16712_1_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_136;
  reg  _T_16712_1_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_137;
  reg  _T_16712_2_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_138;
  reg  _T_16712_2_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_139;
  reg  _T_16712_3_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_140;
  reg  _T_16712_3_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_141;
  reg  _T_16712_4_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_142;
  reg  _T_16712_4_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_143;
  reg  _T_16712_5_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_144;
  reg  _T_16712_5_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_145;
  reg  _T_16712_6_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_146;
  reg  _T_16712_6_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_147;
  reg  _T_16712_7_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_148;
  reg  _T_16712_7_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_149;
  reg  _T_16712_8_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_150;
  reg  _T_16712_8_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_151;
  reg  _T_16712_9_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_152;
  reg  _T_16712_9_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_153;
  reg  _T_16712_10_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_154;
  reg  _T_16712_10_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_155;
  reg  _T_16712_11_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_156;
  reg  _T_16712_11_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_157;
  reg  _T_16712_12_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_158;
  reg  _T_16712_12_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_159;
  reg  _T_16712_13_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_160;
  reg  _T_16712_13_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_161;
  reg  _T_16712_14_0; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_162;
  reg  _T_16712_14_1; // @[Reg.scala 11:16:@2958.4]
  reg [31:0] _RAND_163;
  reg  datRreqd2_0_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_164;
  reg  datRreqd2_0_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_165;
  reg  datRreqd2_1_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_166;
  reg  datRreqd2_1_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_167;
  reg  datRreqd2_2_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_168;
  reg  datRreqd2_2_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_169;
  reg  datRreqd2_3_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_170;
  reg  datRreqd2_3_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_171;
  reg  datRreqd2_4_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_172;
  reg  datRreqd2_4_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_173;
  reg  datRreqd2_5_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_174;
  reg  datRreqd2_5_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_175;
  reg  datRreqd2_6_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_176;
  reg  datRreqd2_6_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_177;
  reg  datRreqd2_7_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_178;
  reg  datRreqd2_7_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_179;
  reg  datRreqd2_8_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_180;
  reg  datRreqd2_8_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_181;
  reg  datRreqd2_9_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_182;
  reg  datRreqd2_9_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_183;
  reg  datRreqd2_10_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_184;
  reg  datRreqd2_10_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_185;
  reg  datRreqd2_11_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_186;
  reg  datRreqd2_11_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_187;
  reg  datRreqd2_12_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_188;
  reg  datRreqd2_12_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_189;
  reg  datRreqd2_13_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_190;
  reg  datRreqd2_13_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_191;
  reg  datRreqd2_14_0; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_192;
  reg  datRreqd2_14_1; // @[Reg.scala 11:16:@2993.4]
  reg [31:0] _RAND_193;
  reg  _T_21752_1_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_194;
  reg  _T_21752_1_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_195;
  reg  _T_21752_2_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_196;
  reg  _T_21752_2_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_197;
  reg  _T_21752_3_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_198;
  reg  _T_21752_3_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_199;
  reg  _T_21752_4_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_200;
  reg  _T_21752_4_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_201;
  reg  _T_21752_5_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_202;
  reg  _T_21752_5_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_203;
  reg  _T_21752_6_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_204;
  reg  _T_21752_6_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_205;
  reg  _T_21752_7_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_206;
  reg  _T_21752_7_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_207;
  reg  _T_21752_8_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_208;
  reg  _T_21752_8_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_209;
  reg  _T_21752_9_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_210;
  reg  _T_21752_9_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_211;
  reg  _T_21752_10_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_212;
  reg  _T_21752_10_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_213;
  reg  _T_21752_11_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_214;
  reg  _T_21752_11_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_215;
  reg  _T_21752_12_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_216;
  reg  _T_21752_12_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_217;
  reg  _T_21752_13_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_218;
  reg  _T_21752_13_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_219;
  reg  _T_21752_14_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_220;
  reg  _T_21752_14_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_221;
  reg  _T_21752_15_0; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_222;
  reg  _T_21752_15_1; // @[Reg.scala 11:16:@3028.4]
  reg [31:0] _RAND_223;
  reg  wtRreqd2_1_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_224;
  reg  wtRreqd2_1_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_225;
  reg  wtRreqd2_2_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_226;
  reg  wtRreqd2_2_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_227;
  reg  wtRreqd2_3_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_228;
  reg  wtRreqd2_3_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_229;
  reg  wtRreqd2_4_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_230;
  reg  wtRreqd2_4_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_231;
  reg  wtRreqd2_5_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_232;
  reg  wtRreqd2_5_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_233;
  reg  wtRreqd2_6_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_234;
  reg  wtRreqd2_6_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_235;
  reg  wtRreqd2_7_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_236;
  reg  wtRreqd2_7_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_237;
  reg  wtRreqd2_8_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_238;
  reg  wtRreqd2_8_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_239;
  reg  wtRreqd2_9_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_240;
  reg  wtRreqd2_9_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_241;
  reg  wtRreqd2_10_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_242;
  reg  wtRreqd2_10_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_243;
  reg  wtRreqd2_11_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_244;
  reg  wtRreqd2_11_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_245;
  reg  wtRreqd2_12_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_246;
  reg  wtRreqd2_12_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_247;
  reg  wtRreqd2_13_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_248;
  reg  wtRreqd2_13_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_249;
  reg  wtRreqd2_14_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_250;
  reg  wtRreqd2_14_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_251;
  reg  wtRreqd2_15_0; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_252;
  reg  wtRreqd2_15_1; // @[Reg.scala 11:16:@3063.4]
  reg [31:0] _RAND_253;
  reg  _T_26101_0; // @[Reg.scala 11:16:@3098.4]
  reg [31:0] _RAND_254;
  reg  _T_26101_1; // @[Reg.scala 11:16:@3098.4]
  reg [31:0] _RAND_255;
  reg  wmbRreqd2_0; // @[Reg.scala 11:16:@3103.4]
  reg [31:0] _RAND_256;
  reg  wmbRreqd2_1; // @[Reg.scala 11:16:@3103.4]
  reg [31:0] _RAND_257;
  reg  _T_26899; // @[Reg.scala 11:16:@3195.4]
  reg [31:0] _RAND_258;
  reg  p0enabled2; // @[Reg.scala 11:16:@3199.4]
  reg [31:0] _RAND_259;
  reg  _T_26903; // @[Reg.scala 11:16:@3203.4]
  reg [31:0] _RAND_260;
  reg  p1enabled2; // @[Reg.scala 11:16:@3207.4]
  reg [31:0] _RAND_261;
  wire [511:0] _T_26912; // @[Bitwise.scala 72:12:@3220.4]
  wire [511:0] _T_26916; // @[Bitwise.scala 72:12:@3222.4]
  wire [1023:0] _T_26917; // @[Cat.scala 30:58:@3223.4]
  wire [511:0] ramdout_0_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3158.4 Cbuf.scala 207:21:@3563.4]
  wire [511:0] ramdout_0_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3157.4 Cbuf.scala 207:21:@3556.4]
  wire [1023:0] _T_26918; // @[Cat.scala 30:58:@3224.4]
  wire [1023:0] _T_26919; // @[Cbuf.scala 186:105:@3225.4]
  wire [511:0] _T_26923; // @[Bitwise.scala 72:12:@3227.4]
  wire [511:0] _T_26927; // @[Bitwise.scala 72:12:@3229.4]
  wire [1023:0] _T_26928; // @[Cat.scala 30:58:@3230.4]
  wire [511:0] ramdout_1_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3160.4 Cbuf.scala 207:21:@3577.4]
  wire [511:0] ramdout_1_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3159.4 Cbuf.scala 207:21:@3570.4]
  wire [1023:0] _T_26929; // @[Cat.scala 30:58:@3231.4]
  wire [1023:0] _T_26930; // @[Cbuf.scala 186:105:@3232.4]
  wire [511:0] _T_26934; // @[Bitwise.scala 72:12:@3234.4]
  wire [511:0] _T_26938; // @[Bitwise.scala 72:12:@3236.4]
  wire [1023:0] _T_26939; // @[Cat.scala 30:58:@3237.4]
  wire [511:0] ramdout_2_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3162.4 Cbuf.scala 207:21:@3591.4]
  wire [511:0] ramdout_2_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3161.4 Cbuf.scala 207:21:@3584.4]
  wire [1023:0] _T_26940; // @[Cat.scala 30:58:@3238.4]
  wire [1023:0] _T_26941; // @[Cbuf.scala 186:105:@3239.4]
  wire [511:0] _T_26945; // @[Bitwise.scala 72:12:@3241.4]
  wire [511:0] _T_26949; // @[Bitwise.scala 72:12:@3243.4]
  wire [1023:0] _T_26950; // @[Cat.scala 30:58:@3244.4]
  wire [511:0] ramdout_3_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3164.4 Cbuf.scala 207:21:@3605.4]
  wire [511:0] ramdout_3_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3163.4 Cbuf.scala 207:21:@3598.4]
  wire [1023:0] _T_26951; // @[Cat.scala 30:58:@3245.4]
  wire [1023:0] _T_26952; // @[Cbuf.scala 186:105:@3246.4]
  wire [511:0] _T_26956; // @[Bitwise.scala 72:12:@3248.4]
  wire [511:0] _T_26960; // @[Bitwise.scala 72:12:@3250.4]
  wire [1023:0] _T_26961; // @[Cat.scala 30:58:@3251.4]
  wire [511:0] ramdout_4_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3166.4 Cbuf.scala 207:21:@3619.4]
  wire [511:0] ramdout_4_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3165.4 Cbuf.scala 207:21:@3612.4]
  wire [1023:0] _T_26962; // @[Cat.scala 30:58:@3252.4]
  wire [1023:0] _T_26963; // @[Cbuf.scala 186:105:@3253.4]
  wire [511:0] _T_26967; // @[Bitwise.scala 72:12:@3255.4]
  wire [511:0] _T_26971; // @[Bitwise.scala 72:12:@3257.4]
  wire [1023:0] _T_26972; // @[Cat.scala 30:58:@3258.4]
  wire [511:0] ramdout_5_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3168.4 Cbuf.scala 207:21:@3633.4]
  wire [511:0] ramdout_5_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3167.4 Cbuf.scala 207:21:@3626.4]
  wire [1023:0] _T_26973; // @[Cat.scala 30:58:@3259.4]
  wire [1023:0] _T_26974; // @[Cbuf.scala 186:105:@3260.4]
  wire [511:0] _T_26978; // @[Bitwise.scala 72:12:@3262.4]
  wire [511:0] _T_26982; // @[Bitwise.scala 72:12:@3264.4]
  wire [1023:0] _T_26983; // @[Cat.scala 30:58:@3265.4]
  wire [511:0] ramdout_6_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3170.4 Cbuf.scala 207:21:@3647.4]
  wire [511:0] ramdout_6_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3169.4 Cbuf.scala 207:21:@3640.4]
  wire [1023:0] _T_26984; // @[Cat.scala 30:58:@3266.4]
  wire [1023:0] _T_26985; // @[Cbuf.scala 186:105:@3267.4]
  wire [511:0] _T_26989; // @[Bitwise.scala 72:12:@3269.4]
  wire [511:0] _T_26993; // @[Bitwise.scala 72:12:@3271.4]
  wire [1023:0] _T_26994; // @[Cat.scala 30:58:@3272.4]
  wire [511:0] ramdout_7_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3172.4 Cbuf.scala 207:21:@3661.4]
  wire [511:0] ramdout_7_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3171.4 Cbuf.scala 207:21:@3654.4]
  wire [1023:0] _T_26995; // @[Cat.scala 30:58:@3273.4]
  wire [1023:0] _T_26996; // @[Cbuf.scala 186:105:@3274.4]
  wire [511:0] _T_27000; // @[Bitwise.scala 72:12:@3276.4]
  wire [511:0] _T_27004; // @[Bitwise.scala 72:12:@3278.4]
  wire [1023:0] _T_27005; // @[Cat.scala 30:58:@3279.4]
  wire [511:0] ramdout_8_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3174.4 Cbuf.scala 207:21:@3675.4]
  wire [511:0] ramdout_8_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3173.4 Cbuf.scala 207:21:@3668.4]
  wire [1023:0] _T_27006; // @[Cat.scala 30:58:@3280.4]
  wire [1023:0] _T_27007; // @[Cbuf.scala 186:105:@3281.4]
  wire [511:0] _T_27011; // @[Bitwise.scala 72:12:@3283.4]
  wire [511:0] _T_27015; // @[Bitwise.scala 72:12:@3285.4]
  wire [1023:0] _T_27016; // @[Cat.scala 30:58:@3286.4]
  wire [511:0] ramdout_9_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3176.4 Cbuf.scala 207:21:@3689.4]
  wire [511:0] ramdout_9_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3175.4 Cbuf.scala 207:21:@3682.4]
  wire [1023:0] _T_27017; // @[Cat.scala 30:58:@3287.4]
  wire [1023:0] _T_27018; // @[Cbuf.scala 186:105:@3288.4]
  wire [511:0] _T_27022; // @[Bitwise.scala 72:12:@3290.4]
  wire [511:0] _T_27026; // @[Bitwise.scala 72:12:@3292.4]
  wire [1023:0] _T_27027; // @[Cat.scala 30:58:@3293.4]
  wire [511:0] ramdout_10_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3178.4 Cbuf.scala 207:21:@3703.4]
  wire [511:0] ramdout_10_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3177.4 Cbuf.scala 207:21:@3696.4]
  wire [1023:0] _T_27028; // @[Cat.scala 30:58:@3294.4]
  wire [1023:0] _T_27029; // @[Cbuf.scala 186:105:@3295.4]
  wire [511:0] _T_27033; // @[Bitwise.scala 72:12:@3297.4]
  wire [511:0] _T_27037; // @[Bitwise.scala 72:12:@3299.4]
  wire [1023:0] _T_27038; // @[Cat.scala 30:58:@3300.4]
  wire [511:0] ramdout_11_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3180.4 Cbuf.scala 207:21:@3717.4]
  wire [511:0] ramdout_11_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3179.4 Cbuf.scala 207:21:@3710.4]
  wire [1023:0] _T_27039; // @[Cat.scala 30:58:@3301.4]
  wire [1023:0] _T_27040; // @[Cbuf.scala 186:105:@3302.4]
  wire [511:0] _T_27044; // @[Bitwise.scala 72:12:@3304.4]
  wire [511:0] _T_27048; // @[Bitwise.scala 72:12:@3306.4]
  wire [1023:0] _T_27049; // @[Cat.scala 30:58:@3307.4]
  wire [511:0] ramdout_12_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3182.4 Cbuf.scala 207:21:@3731.4]
  wire [511:0] ramdout_12_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3181.4 Cbuf.scala 207:21:@3724.4]
  wire [1023:0] _T_27050; // @[Cat.scala 30:58:@3308.4]
  wire [1023:0] _T_27051; // @[Cbuf.scala 186:105:@3309.4]
  wire [511:0] _T_27055; // @[Bitwise.scala 72:12:@3311.4]
  wire [511:0] _T_27059; // @[Bitwise.scala 72:12:@3313.4]
  wire [1023:0] _T_27060; // @[Cat.scala 30:58:@3314.4]
  wire [511:0] ramdout_13_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3184.4 Cbuf.scala 207:21:@3745.4]
  wire [511:0] ramdout_13_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3183.4 Cbuf.scala 207:21:@3738.4]
  wire [1023:0] _T_27061; // @[Cat.scala 30:58:@3315.4]
  wire [1023:0] _T_27062; // @[Cbuf.scala 186:105:@3316.4]
  wire [511:0] _T_27066; // @[Bitwise.scala 72:12:@3318.4]
  wire [511:0] _T_27070; // @[Bitwise.scala 72:12:@3320.4]
  wire [1023:0] _T_27071; // @[Cat.scala 30:58:@3321.4]
  wire [511:0] ramdout_14_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3186.4 Cbuf.scala 207:21:@3759.4]
  wire [511:0] ramdout_14_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3185.4 Cbuf.scala 207:21:@3752.4]
  wire [1023:0] _T_27072; // @[Cat.scala 30:58:@3322.4]
  wire [1023:0] _T_27073; // @[Cbuf.scala 186:105:@3323.4]
  wire [1023:0] _T_27074; // @[Cbuf.scala 186:151:@3324.4]
  wire [1023:0] _T_27075; // @[Cbuf.scala 186:151:@3325.4]
  wire [1023:0] _T_27076; // @[Cbuf.scala 186:151:@3326.4]
  wire [1023:0] _T_27077; // @[Cbuf.scala 186:151:@3327.4]
  wire [1023:0] _T_27078; // @[Cbuf.scala 186:151:@3328.4]
  wire [1023:0] _T_27079; // @[Cbuf.scala 186:151:@3329.4]
  wire [1023:0] _T_27080; // @[Cbuf.scala 186:151:@3330.4]
  wire [1023:0] _T_27081; // @[Cbuf.scala 186:151:@3331.4]
  wire [1023:0] _T_27082; // @[Cbuf.scala 186:151:@3332.4]
  wire [1023:0] _T_27083; // @[Cbuf.scala 186:151:@3333.4]
  wire [1023:0] _T_27084; // @[Cbuf.scala 186:151:@3334.4]
  wire [1023:0] _T_27085; // @[Cbuf.scala 186:151:@3335.4]
  wire [1023:0] _T_27086; // @[Cbuf.scala 186:151:@3336.4]
  reg [1023:0] p0Datad3; // @[Cbuf.scala 186:22:@3338.4]
  reg [1023:0] _RAND_262;
  reg  p0Validd3; // @[Cbuf.scala 187:23:@3341.4]
  reg [31:0] _RAND_263;
  wire [511:0] _T_27095; // @[Bitwise.scala 72:12:@3345.4]
  wire [511:0] _T_27099; // @[Bitwise.scala 72:12:@3347.4]
  wire [1023:0] _T_27100; // @[Cat.scala 30:58:@3348.4]
  wire [1023:0] _T_27102; // @[Cbuf.scala 188:103:@3350.4]
  wire [511:0] _T_27106; // @[Bitwise.scala 72:12:@3352.4]
  wire [511:0] _T_27110; // @[Bitwise.scala 72:12:@3354.4]
  wire [1023:0] _T_27111; // @[Cat.scala 30:58:@3355.4]
  wire [1023:0] _T_27113; // @[Cbuf.scala 188:103:@3357.4]
  wire [511:0] _T_27117; // @[Bitwise.scala 72:12:@3359.4]
  wire [511:0] _T_27121; // @[Bitwise.scala 72:12:@3361.4]
  wire [1023:0] _T_27122; // @[Cat.scala 30:58:@3362.4]
  wire [1023:0] _T_27124; // @[Cbuf.scala 188:103:@3364.4]
  wire [511:0] _T_27128; // @[Bitwise.scala 72:12:@3366.4]
  wire [511:0] _T_27132; // @[Bitwise.scala 72:12:@3368.4]
  wire [1023:0] _T_27133; // @[Cat.scala 30:58:@3369.4]
  wire [1023:0] _T_27135; // @[Cbuf.scala 188:103:@3371.4]
  wire [511:0] _T_27139; // @[Bitwise.scala 72:12:@3373.4]
  wire [511:0] _T_27143; // @[Bitwise.scala 72:12:@3375.4]
  wire [1023:0] _T_27144; // @[Cat.scala 30:58:@3376.4]
  wire [1023:0] _T_27146; // @[Cbuf.scala 188:103:@3378.4]
  wire [511:0] _T_27150; // @[Bitwise.scala 72:12:@3380.4]
  wire [511:0] _T_27154; // @[Bitwise.scala 72:12:@3382.4]
  wire [1023:0] _T_27155; // @[Cat.scala 30:58:@3383.4]
  wire [1023:0] _T_27157; // @[Cbuf.scala 188:103:@3385.4]
  wire [511:0] _T_27161; // @[Bitwise.scala 72:12:@3387.4]
  wire [511:0] _T_27165; // @[Bitwise.scala 72:12:@3389.4]
  wire [1023:0] _T_27166; // @[Cat.scala 30:58:@3390.4]
  wire [1023:0] _T_27168; // @[Cbuf.scala 188:103:@3392.4]
  wire [511:0] _T_27172; // @[Bitwise.scala 72:12:@3394.4]
  wire [511:0] _T_27176; // @[Bitwise.scala 72:12:@3396.4]
  wire [1023:0] _T_27177; // @[Cat.scala 30:58:@3397.4]
  wire [1023:0] _T_27179; // @[Cbuf.scala 188:103:@3399.4]
  wire [511:0] _T_27183; // @[Bitwise.scala 72:12:@3401.4]
  wire [511:0] _T_27187; // @[Bitwise.scala 72:12:@3403.4]
  wire [1023:0] _T_27188; // @[Cat.scala 30:58:@3404.4]
  wire [1023:0] _T_27190; // @[Cbuf.scala 188:103:@3406.4]
  wire [511:0] _T_27194; // @[Bitwise.scala 72:12:@3408.4]
  wire [511:0] _T_27198; // @[Bitwise.scala 72:12:@3410.4]
  wire [1023:0] _T_27199; // @[Cat.scala 30:58:@3411.4]
  wire [1023:0] _T_27201; // @[Cbuf.scala 188:103:@3413.4]
  wire [511:0] _T_27205; // @[Bitwise.scala 72:12:@3415.4]
  wire [511:0] _T_27209; // @[Bitwise.scala 72:12:@3417.4]
  wire [1023:0] _T_27210; // @[Cat.scala 30:58:@3418.4]
  wire [1023:0] _T_27212; // @[Cbuf.scala 188:103:@3420.4]
  wire [511:0] _T_27216; // @[Bitwise.scala 72:12:@3422.4]
  wire [511:0] _T_27220; // @[Bitwise.scala 72:12:@3424.4]
  wire [1023:0] _T_27221; // @[Cat.scala 30:58:@3425.4]
  wire [1023:0] _T_27223; // @[Cbuf.scala 188:103:@3427.4]
  wire [511:0] _T_27227; // @[Bitwise.scala 72:12:@3429.4]
  wire [511:0] _T_27231; // @[Bitwise.scala 72:12:@3431.4]
  wire [1023:0] _T_27232; // @[Cat.scala 30:58:@3432.4]
  wire [1023:0] _T_27234; // @[Cbuf.scala 188:103:@3434.4]
  wire [511:0] _T_27238; // @[Bitwise.scala 72:12:@3436.4]
  wire [511:0] _T_27242; // @[Bitwise.scala 72:12:@3438.4]
  wire [1023:0] _T_27243; // @[Cat.scala 30:58:@3439.4]
  wire [1023:0] _T_27245; // @[Cbuf.scala 188:103:@3441.4]
  wire [511:0] _T_27249; // @[Bitwise.scala 72:12:@3443.4]
  wire [511:0] _T_27253; // @[Bitwise.scala 72:12:@3445.4]
  wire [1023:0] _T_27254; // @[Cat.scala 30:58:@3446.4]
  wire [511:0] ramdout_15_1; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3188.4 Cbuf.scala 207:21:@3773.4]
  wire [511:0] ramdout_15_0; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3187.4 Cbuf.scala 207:21:@3766.4]
  wire [1023:0] _T_27255; // @[Cat.scala 30:58:@3447.4]
  wire [1023:0] _T_27256; // @[Cbuf.scala 188:103:@3448.4]
  wire [1023:0] _T_27257; // @[Cbuf.scala 188:149:@3449.4]
  wire [1023:0] _T_27258; // @[Cbuf.scala 188:149:@3450.4]
  wire [1023:0] _T_27259; // @[Cbuf.scala 188:149:@3451.4]
  wire [1023:0] _T_27260; // @[Cbuf.scala 188:149:@3452.4]
  wire [1023:0] _T_27261; // @[Cbuf.scala 188:149:@3453.4]
  wire [1023:0] _T_27262; // @[Cbuf.scala 188:149:@3454.4]
  wire [1023:0] _T_27263; // @[Cbuf.scala 188:149:@3455.4]
  wire [1023:0] _T_27264; // @[Cbuf.scala 188:149:@3456.4]
  wire [1023:0] _T_27265; // @[Cbuf.scala 188:149:@3457.4]
  wire [1023:0] _T_27266; // @[Cbuf.scala 188:149:@3458.4]
  wire [1023:0] _T_27267; // @[Cbuf.scala 188:149:@3459.4]
  wire [1023:0] _T_27268; // @[Cbuf.scala 188:149:@3460.4]
  wire [1023:0] _T_27269; // @[Cbuf.scala 188:149:@3461.4]
  reg [1023:0] p1Datad3; // @[Cbuf.scala 188:22:@3463.4]
  reg [1023:0] _RAND_264;
  reg  p1Validd3; // @[Cbuf.scala 189:23:@3466.4]
  reg [31:0] _RAND_265;
  wire [511:0] _T_27278; // @[Bitwise.scala 72:12:@3470.4]
  wire [511:0] _T_27282; // @[Bitwise.scala 72:12:@3472.4]
  wire [1023:0] _T_27283; // @[Cat.scala 30:58:@3473.4]
  reg [1023:0] p2Datad3; // @[Cbuf.scala 190:22:@3476.4]
  reg [1023:0] _RAND_266;
  reg  p2Validd3; // @[Cbuf.scala 191:23:@3479.4]
  reg [31:0] _RAND_267;
  reg [1023:0] _T_27292; // @[Reg.scala 11:16:@3482.4]
  reg [1023:0] _RAND_268;
  reg [1023:0] _T_27294; // @[Reg.scala 11:16:@3486.4]
  reg [1023:0] _RAND_269;
  reg [1023:0] p0Datad6; // @[Reg.scala 11:16:@3490.4]
  reg [1023:0] _RAND_270;
  reg  _T_27298; // @[Reg.scala 11:16:@3494.4]
  reg [31:0] _RAND_271;
  reg  _T_27300; // @[Reg.scala 11:16:@3498.4]
  reg [31:0] _RAND_272;
  reg  p0Validd6; // @[Reg.scala 11:16:@3502.4]
  reg [31:0] _RAND_273;
  reg [1023:0] _T_27304; // @[Reg.scala 11:16:@3506.4]
  reg [1023:0] _RAND_274;
  reg [1023:0] _T_27306; // @[Reg.scala 11:16:@3510.4]
  reg [1023:0] _RAND_275;
  reg [1023:0] p1Datad6; // @[Reg.scala 11:16:@3514.4]
  reg [1023:0] _RAND_276;
  reg  _T_27310; // @[Reg.scala 11:16:@3518.4]
  reg [31:0] _RAND_277;
  reg  _T_27312; // @[Reg.scala 11:16:@3522.4]
  reg [31:0] _RAND_278;
  reg  p1Validd6; // @[Reg.scala 11:16:@3526.4]
  reg [31:0] _RAND_279;
  reg [1023:0] _T_27316; // @[Reg.scala 11:16:@3530.4]
  reg [1023:0] _RAND_280;
  reg [1023:0] _T_27318; // @[Reg.scala 11:16:@3534.4]
  reg [1023:0] _RAND_281;
  reg [1023:0] p2Datad6; // @[Reg.scala 11:16:@3538.4]
  reg [1023:0] _RAND_282;
  reg  _T_27322; // @[Reg.scala 11:16:@3542.4]
  reg [31:0] _RAND_283;
  reg  _T_27324; // @[Reg.scala 11:16:@3546.4]
  reg [31:0] _RAND_284;
  reg  p2Validd6; // @[Reg.scala 11:16:@3550.4]
  reg [31:0] _RAND_285;
  RamSync RamSync ( // @[Cbuf.scala 43:52:@648.4]
    .clock(RamSync_clock),
    .io_re(RamSync_io_re),
    .io_we(RamSync_io_we),
    .io_ra(RamSync_io_ra),
    .io_wa(RamSync_io_wa),
    .io_di(RamSync_io_di),
    .io_dout(RamSync_io_dout)
  );
  RamSync RamSync_1 ( // @[Cbuf.scala 43:52:@651.4]
    .clock(RamSync_1_clock),
    .io_re(RamSync_1_io_re),
    .io_we(RamSync_1_io_we),
    .io_ra(RamSync_1_io_ra),
    .io_wa(RamSync_1_io_wa),
    .io_di(RamSync_1_io_di),
    .io_dout(RamSync_1_io_dout)
  );
  RamSync RamSync_2 ( // @[Cbuf.scala 43:52:@654.4]
    .clock(RamSync_2_clock),
    .io_re(RamSync_2_io_re),
    .io_we(RamSync_2_io_we),
    .io_ra(RamSync_2_io_ra),
    .io_wa(RamSync_2_io_wa),
    .io_di(RamSync_2_io_di),
    .io_dout(RamSync_2_io_dout)
  );
  RamSync RamSync_3 ( // @[Cbuf.scala 43:52:@657.4]
    .clock(RamSync_3_clock),
    .io_re(RamSync_3_io_re),
    .io_we(RamSync_3_io_we),
    .io_ra(RamSync_3_io_ra),
    .io_wa(RamSync_3_io_wa),
    .io_di(RamSync_3_io_di),
    .io_dout(RamSync_3_io_dout)
  );
  RamSync RamSync_4 ( // @[Cbuf.scala 43:52:@660.4]
    .clock(RamSync_4_clock),
    .io_re(RamSync_4_io_re),
    .io_we(RamSync_4_io_we),
    .io_ra(RamSync_4_io_ra),
    .io_wa(RamSync_4_io_wa),
    .io_di(RamSync_4_io_di),
    .io_dout(RamSync_4_io_dout)
  );
  RamSync RamSync_5 ( // @[Cbuf.scala 43:52:@663.4]
    .clock(RamSync_5_clock),
    .io_re(RamSync_5_io_re),
    .io_we(RamSync_5_io_we),
    .io_ra(RamSync_5_io_ra),
    .io_wa(RamSync_5_io_wa),
    .io_di(RamSync_5_io_di),
    .io_dout(RamSync_5_io_dout)
  );
  RamSync RamSync_6 ( // @[Cbuf.scala 43:52:@666.4]
    .clock(RamSync_6_clock),
    .io_re(RamSync_6_io_re),
    .io_we(RamSync_6_io_we),
    .io_ra(RamSync_6_io_ra),
    .io_wa(RamSync_6_io_wa),
    .io_di(RamSync_6_io_di),
    .io_dout(RamSync_6_io_dout)
  );
  RamSync RamSync_7 ( // @[Cbuf.scala 43:52:@669.4]
    .clock(RamSync_7_clock),
    .io_re(RamSync_7_io_re),
    .io_we(RamSync_7_io_we),
    .io_ra(RamSync_7_io_ra),
    .io_wa(RamSync_7_io_wa),
    .io_di(RamSync_7_io_di),
    .io_dout(RamSync_7_io_dout)
  );
  RamSync RamSync_8 ( // @[Cbuf.scala 43:52:@672.4]
    .clock(RamSync_8_clock),
    .io_re(RamSync_8_io_re),
    .io_we(RamSync_8_io_we),
    .io_ra(RamSync_8_io_ra),
    .io_wa(RamSync_8_io_wa),
    .io_di(RamSync_8_io_di),
    .io_dout(RamSync_8_io_dout)
  );
  RamSync RamSync_9 ( // @[Cbuf.scala 43:52:@675.4]
    .clock(RamSync_9_clock),
    .io_re(RamSync_9_io_re),
    .io_we(RamSync_9_io_we),
    .io_ra(RamSync_9_io_ra),
    .io_wa(RamSync_9_io_wa),
    .io_di(RamSync_9_io_di),
    .io_dout(RamSync_9_io_dout)
  );
  RamSync RamSync_10 ( // @[Cbuf.scala 43:52:@678.4]
    .clock(RamSync_10_clock),
    .io_re(RamSync_10_io_re),
    .io_we(RamSync_10_io_we),
    .io_ra(RamSync_10_io_ra),
    .io_wa(RamSync_10_io_wa),
    .io_di(RamSync_10_io_di),
    .io_dout(RamSync_10_io_dout)
  );
  RamSync RamSync_11 ( // @[Cbuf.scala 43:52:@681.4]
    .clock(RamSync_11_clock),
    .io_re(RamSync_11_io_re),
    .io_we(RamSync_11_io_we),
    .io_ra(RamSync_11_io_ra),
    .io_wa(RamSync_11_io_wa),
    .io_di(RamSync_11_io_di),
    .io_dout(RamSync_11_io_dout)
  );
  RamSync RamSync_12 ( // @[Cbuf.scala 43:52:@684.4]
    .clock(RamSync_12_clock),
    .io_re(RamSync_12_io_re),
    .io_we(RamSync_12_io_we),
    .io_ra(RamSync_12_io_ra),
    .io_wa(RamSync_12_io_wa),
    .io_di(RamSync_12_io_di),
    .io_dout(RamSync_12_io_dout)
  );
  RamSync RamSync_13 ( // @[Cbuf.scala 43:52:@687.4]
    .clock(RamSync_13_clock),
    .io_re(RamSync_13_io_re),
    .io_we(RamSync_13_io_we),
    .io_ra(RamSync_13_io_ra),
    .io_wa(RamSync_13_io_wa),
    .io_di(RamSync_13_io_di),
    .io_dout(RamSync_13_io_dout)
  );
  RamSync RamSync_14 ( // @[Cbuf.scala 43:52:@690.4]
    .clock(RamSync_14_clock),
    .io_re(RamSync_14_io_re),
    .io_we(RamSync_14_io_we),
    .io_ra(RamSync_14_io_ra),
    .io_wa(RamSync_14_io_wa),
    .io_di(RamSync_14_io_di),
    .io_dout(RamSync_14_io_dout)
  );
  RamSync RamSync_15 ( // @[Cbuf.scala 43:52:@693.4]
    .clock(RamSync_15_clock),
    .io_re(RamSync_15_io_re),
    .io_we(RamSync_15_io_we),
    .io_ra(RamSync_15_io_ra),
    .io_wa(RamSync_15_io_wa),
    .io_di(RamSync_15_io_di),
    .io_dout(RamSync_15_io_dout)
  );
  RamSync RamSync_16 ( // @[Cbuf.scala 43:52:@696.4]
    .clock(RamSync_16_clock),
    .io_re(RamSync_16_io_re),
    .io_we(RamSync_16_io_we),
    .io_ra(RamSync_16_io_ra),
    .io_wa(RamSync_16_io_wa),
    .io_di(RamSync_16_io_di),
    .io_dout(RamSync_16_io_dout)
  );
  RamSync RamSync_17 ( // @[Cbuf.scala 43:52:@699.4]
    .clock(RamSync_17_clock),
    .io_re(RamSync_17_io_re),
    .io_we(RamSync_17_io_we),
    .io_ra(RamSync_17_io_ra),
    .io_wa(RamSync_17_io_wa),
    .io_di(RamSync_17_io_di),
    .io_dout(RamSync_17_io_dout)
  );
  RamSync RamSync_18 ( // @[Cbuf.scala 43:52:@702.4]
    .clock(RamSync_18_clock),
    .io_re(RamSync_18_io_re),
    .io_we(RamSync_18_io_we),
    .io_ra(RamSync_18_io_ra),
    .io_wa(RamSync_18_io_wa),
    .io_di(RamSync_18_io_di),
    .io_dout(RamSync_18_io_dout)
  );
  RamSync RamSync_19 ( // @[Cbuf.scala 43:52:@705.4]
    .clock(RamSync_19_clock),
    .io_re(RamSync_19_io_re),
    .io_we(RamSync_19_io_we),
    .io_ra(RamSync_19_io_ra),
    .io_wa(RamSync_19_io_wa),
    .io_di(RamSync_19_io_di),
    .io_dout(RamSync_19_io_dout)
  );
  RamSync RamSync_20 ( // @[Cbuf.scala 43:52:@708.4]
    .clock(RamSync_20_clock),
    .io_re(RamSync_20_io_re),
    .io_we(RamSync_20_io_we),
    .io_ra(RamSync_20_io_ra),
    .io_wa(RamSync_20_io_wa),
    .io_di(RamSync_20_io_di),
    .io_dout(RamSync_20_io_dout)
  );
  RamSync RamSync_21 ( // @[Cbuf.scala 43:52:@711.4]
    .clock(RamSync_21_clock),
    .io_re(RamSync_21_io_re),
    .io_we(RamSync_21_io_we),
    .io_ra(RamSync_21_io_ra),
    .io_wa(RamSync_21_io_wa),
    .io_di(RamSync_21_io_di),
    .io_dout(RamSync_21_io_dout)
  );
  RamSync RamSync_22 ( // @[Cbuf.scala 43:52:@714.4]
    .clock(RamSync_22_clock),
    .io_re(RamSync_22_io_re),
    .io_we(RamSync_22_io_we),
    .io_ra(RamSync_22_io_ra),
    .io_wa(RamSync_22_io_wa),
    .io_di(RamSync_22_io_di),
    .io_dout(RamSync_22_io_dout)
  );
  RamSync RamSync_23 ( // @[Cbuf.scala 43:52:@717.4]
    .clock(RamSync_23_clock),
    .io_re(RamSync_23_io_re),
    .io_we(RamSync_23_io_we),
    .io_ra(RamSync_23_io_ra),
    .io_wa(RamSync_23_io_wa),
    .io_di(RamSync_23_io_di),
    .io_dout(RamSync_23_io_dout)
  );
  RamSync RamSync_24 ( // @[Cbuf.scala 43:52:@720.4]
    .clock(RamSync_24_clock),
    .io_re(RamSync_24_io_re),
    .io_we(RamSync_24_io_we),
    .io_ra(RamSync_24_io_ra),
    .io_wa(RamSync_24_io_wa),
    .io_di(RamSync_24_io_di),
    .io_dout(RamSync_24_io_dout)
  );
  RamSync RamSync_25 ( // @[Cbuf.scala 43:52:@723.4]
    .clock(RamSync_25_clock),
    .io_re(RamSync_25_io_re),
    .io_we(RamSync_25_io_we),
    .io_ra(RamSync_25_io_ra),
    .io_wa(RamSync_25_io_wa),
    .io_di(RamSync_25_io_di),
    .io_dout(RamSync_25_io_dout)
  );
  RamSync RamSync_26 ( // @[Cbuf.scala 43:52:@726.4]
    .clock(RamSync_26_clock),
    .io_re(RamSync_26_io_re),
    .io_we(RamSync_26_io_we),
    .io_ra(RamSync_26_io_ra),
    .io_wa(RamSync_26_io_wa),
    .io_di(RamSync_26_io_di),
    .io_dout(RamSync_26_io_dout)
  );
  RamSync RamSync_27 ( // @[Cbuf.scala 43:52:@729.4]
    .clock(RamSync_27_clock),
    .io_re(RamSync_27_io_re),
    .io_we(RamSync_27_io_we),
    .io_ra(RamSync_27_io_ra),
    .io_wa(RamSync_27_io_wa),
    .io_di(RamSync_27_io_di),
    .io_dout(RamSync_27_io_dout)
  );
  RamSync RamSync_28 ( // @[Cbuf.scala 43:52:@732.4]
    .clock(RamSync_28_clock),
    .io_re(RamSync_28_io_re),
    .io_we(RamSync_28_io_we),
    .io_ra(RamSync_28_io_ra),
    .io_wa(RamSync_28_io_wa),
    .io_di(RamSync_28_io_di),
    .io_dout(RamSync_28_io_dout)
  );
  RamSync RamSync_29 ( // @[Cbuf.scala 43:52:@735.4]
    .clock(RamSync_29_clock),
    .io_re(RamSync_29_io_re),
    .io_we(RamSync_29_io_we),
    .io_ra(RamSync_29_io_ra),
    .io_wa(RamSync_29_io_wa),
    .io_di(RamSync_29_io_di),
    .io_dout(RamSync_29_io_dout)
  );
  RamSync RamSync_30 ( // @[Cbuf.scala 43:52:@738.4]
    .clock(RamSync_30_clock),
    .io_re(RamSync_30_io_re),
    .io_we(RamSync_30_io_we),
    .io_ra(RamSync_30_io_ra),
    .io_wa(RamSync_30_io_wa),
    .io_di(RamSync_30_io_di),
    .io_dout(RamSync_30_io_dout)
  );
  RamSync RamSync_31 ( // @[Cbuf.scala 43:52:@741.4]
    .clock(RamSync_31_clock),
    .io_re(RamSync_31_io_re),
    .io_we(RamSync_31_io_we),
    .io_ra(RamSync_31_io_ra),
    .io_wa(RamSync_31_io_wa),
    .io_di(RamSync_31_io_di),
    .io_dout(RamSync_31_io_dout)
  );
  assign _T_1533 = io_cdma2bufDat_addr[11:8]; // @[Cbuf.scala 54:30:@906.4]
  assign _T_1558 = io_cdma2bufDat_hsel[0]; // @[Cbuf.scala 54:87:@907.4]
  assign _T_1559 = io_cdma2bufDat_enable & _T_1558; // @[Cbuf.scala 54:66:@908.4]
  assign datWreq_0_0 = 4'h0 == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_1_0 = 4'h1 == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_2_0 = 4'h2 == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_3_0 = 4'h3 == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_4_0 = 4'h4 == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_5_0 = 4'h5 == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_6_0 = 4'h6 == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_7_0 = 4'h7 == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_8_0 = 4'h8 == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_9_0 = 4'h9 == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_10_0 = 4'ha == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_11_0 = 4'hb == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_12_0 = 4'hc == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_13_0 = 4'hd == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign datWreq_14_0 = 4'he == _T_1533 ? _T_1559 : 1'h0; // @[Cbuf.scala 54:41:@909.4]
  assign _T_1585 = io_cdma2bufDat_hsel[1]; // @[Cbuf.scala 55:87:@911.4]
  assign _T_1586 = io_cdma2bufDat_enable & _T_1585; // @[Cbuf.scala 55:66:@912.4]
  assign datWreq_0_1 = 4'h0 == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_1_1 = 4'h1 == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_2_1 = 4'h2 == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_3_1 = 4'h3 == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_4_1 = 4'h4 == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_5_1 = 4'h5 == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_6_1 = 4'h6 == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_7_1 = 4'h7 == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_8_1 = 4'h8 == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_9_1 = 4'h9 == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_10_1 = 4'ha == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_11_1 = 4'hb == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_12_1 = 4'hc == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_13_1 = 4'hd == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign datWreq_14_1 = 4'he == _T_1533 ? _T_1586 : 1'h0; // @[Cbuf.scala 55:41:@913.4]
  assign _T_1587 = io_cdma2bufWt_addr[11:8]; // @[Cbuf.scala 58:28:@914.4]
  assign _T_1612 = io_cdma2bufWt_hsel[0]; // @[Cbuf.scala 58:85:@915.4]
  assign _T_1614 = _T_1612 == 1'h0; // @[Cbuf.scala 58:66:@916.4]
  assign _T_1615 = io_cdma2bufWt_enable & _T_1614; // @[Cbuf.scala 58:63:@917.4]
  assign wtWreq_1_0 = 4'h1 == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_2_0 = 4'h2 == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_3_0 = 4'h3 == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_4_0 = 4'h4 == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_5_0 = 4'h5 == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_6_0 = 4'h6 == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_7_0 = 4'h7 == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_8_0 = 4'h8 == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_9_0 = 4'h9 == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_10_0 = 4'ha == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_11_0 = 4'hb == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_12_0 = 4'hc == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_13_0 = 4'hd == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_14_0 = 4'he == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign wtWreq_15_0 = 4'hf == _T_1587 ? _T_1615 : 1'h0; // @[Cbuf.scala 58:39:@918.4]
  assign _T_1642 = io_cdma2bufWt_enable & _T_1612; // @[Cbuf.scala 59:63:@921.4]
  assign wtWreq_1_1 = 4'h1 == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_2_1 = 4'h2 == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_3_1 = 4'h3 == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_4_1 = 4'h4 == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_5_1 = 4'h5 == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_6_1 = 4'h6 == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_7_1 = 4'h7 == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_8_1 = 4'h8 == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_9_1 = 4'h9 == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_10_1 = 4'ha == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_11_1 = 4'hb == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_12_1 = 4'hc == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_13_1 = 4'hd == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_14_1 = 4'he == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign wtWreq_15_1 = 4'hf == _T_1587 ? _T_1642 : 1'h0; // @[Cbuf.scala 59:39:@922.4]
  assign _T_4142 = datWreq_1_0 | wtWreq_1_0; // @[Cbuf.scala 84:40:@1025.4]
  assign _T_4143 = datWreq_1_1 | wtWreq_1_1; // @[Cbuf.scala 85:40:@1027.4]
  assign _T_4144 = datWreq_2_0 | wtWreq_2_0; // @[Cbuf.scala 84:40:@1029.4]
  assign _T_4145 = datWreq_2_1 | wtWreq_2_1; // @[Cbuf.scala 85:40:@1031.4]
  assign _T_4146 = datWreq_3_0 | wtWreq_3_0; // @[Cbuf.scala 84:40:@1033.4]
  assign _T_4147 = datWreq_3_1 | wtWreq_3_1; // @[Cbuf.scala 85:40:@1035.4]
  assign _T_4148 = datWreq_4_0 | wtWreq_4_0; // @[Cbuf.scala 84:40:@1037.4]
  assign _T_4149 = datWreq_4_1 | wtWreq_4_1; // @[Cbuf.scala 85:40:@1039.4]
  assign _T_4150 = datWreq_5_0 | wtWreq_5_0; // @[Cbuf.scala 84:40:@1041.4]
  assign _T_4151 = datWreq_5_1 | wtWreq_5_1; // @[Cbuf.scala 85:40:@1043.4]
  assign _T_4152 = datWreq_6_0 | wtWreq_6_0; // @[Cbuf.scala 84:40:@1045.4]
  assign _T_4153 = datWreq_6_1 | wtWreq_6_1; // @[Cbuf.scala 85:40:@1047.4]
  assign _T_4154 = datWreq_7_0 | wtWreq_7_0; // @[Cbuf.scala 84:40:@1049.4]
  assign _T_4155 = datWreq_7_1 | wtWreq_7_1; // @[Cbuf.scala 85:40:@1051.4]
  assign _T_4156 = datWreq_8_0 | wtWreq_8_0; // @[Cbuf.scala 84:40:@1053.4]
  assign _T_4157 = datWreq_8_1 | wtWreq_8_1; // @[Cbuf.scala 85:40:@1055.4]
  assign _T_4158 = datWreq_9_0 | wtWreq_9_0; // @[Cbuf.scala 84:40:@1057.4]
  assign _T_4159 = datWreq_9_1 | wtWreq_9_1; // @[Cbuf.scala 85:40:@1059.4]
  assign _T_4160 = datWreq_10_0 | wtWreq_10_0; // @[Cbuf.scala 84:40:@1061.4]
  assign _T_4161 = datWreq_10_1 | wtWreq_10_1; // @[Cbuf.scala 85:40:@1063.4]
  assign _T_4162 = datWreq_11_0 | wtWreq_11_0; // @[Cbuf.scala 84:40:@1065.4]
  assign _T_4163 = datWreq_11_1 | wtWreq_11_1; // @[Cbuf.scala 85:40:@1067.4]
  assign _T_4164 = datWreq_12_0 | wtWreq_12_0; // @[Cbuf.scala 84:40:@1069.4]
  assign _T_4165 = datWreq_12_1 | wtWreq_12_1; // @[Cbuf.scala 85:40:@1071.4]
  assign _T_4166 = datWreq_13_0 | wtWreq_13_0; // @[Cbuf.scala 84:40:@1073.4]
  assign _T_4167 = datWreq_13_1 | wtWreq_13_1; // @[Cbuf.scala 85:40:@1075.4]
  assign _T_4168 = datWreq_14_0 | wtWreq_14_0; // @[Cbuf.scala 84:40:@1077.4]
  assign _T_4169 = datWreq_14_1 | wtWreq_14_1; // @[Cbuf.scala 85:40:@1079.4]
  assign _T_5162 = ramWreqd1_1_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1465.4]
  assign _T_5166 = ramWreqd1_1_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1467.4]
  assign _T_5171 = ramWreqd1_1_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1471.4]
  assign _T_5175 = ramWreqd1_1_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1473.4]
  assign _T_5180 = ramWreqd1_1_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1477.4]
  assign _T_5184 = ramWreqd1_1_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1479.4]
  assign _T_5189 = ramWreqd1_1_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1483.4]
  assign _T_5193 = ramWreqd1_1_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1485.4]
  assign _T_5198 = ramWreqd1_2_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1489.4]
  assign _T_5202 = ramWreqd1_2_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1491.4]
  assign _T_5207 = ramWreqd1_2_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1495.4]
  assign _T_5211 = ramWreqd1_2_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1497.4]
  assign _T_5216 = ramWreqd1_2_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1501.4]
  assign _T_5220 = ramWreqd1_2_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1503.4]
  assign _T_5225 = ramWreqd1_2_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1507.4]
  assign _T_5229 = ramWreqd1_2_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1509.4]
  assign _T_5234 = ramWreqd1_3_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1513.4]
  assign _T_5238 = ramWreqd1_3_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1515.4]
  assign _T_5243 = ramWreqd1_3_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1519.4]
  assign _T_5247 = ramWreqd1_3_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1521.4]
  assign _T_5252 = ramWreqd1_3_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1525.4]
  assign _T_5256 = ramWreqd1_3_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1527.4]
  assign _T_5261 = ramWreqd1_3_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1531.4]
  assign _T_5265 = ramWreqd1_3_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1533.4]
  assign _T_5270 = ramWreqd1_4_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1537.4]
  assign _T_5274 = ramWreqd1_4_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1539.4]
  assign _T_5279 = ramWreqd1_4_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1543.4]
  assign _T_5283 = ramWreqd1_4_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1545.4]
  assign _T_5288 = ramWreqd1_4_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1549.4]
  assign _T_5292 = ramWreqd1_4_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1551.4]
  assign _T_5297 = ramWreqd1_4_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1555.4]
  assign _T_5301 = ramWreqd1_4_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1557.4]
  assign _T_5306 = ramWreqd1_5_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1561.4]
  assign _T_5310 = ramWreqd1_5_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1563.4]
  assign _T_5315 = ramWreqd1_5_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1567.4]
  assign _T_5319 = ramWreqd1_5_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1569.4]
  assign _T_5324 = ramWreqd1_5_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1573.4]
  assign _T_5328 = ramWreqd1_5_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1575.4]
  assign _T_5333 = ramWreqd1_5_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1579.4]
  assign _T_5337 = ramWreqd1_5_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1581.4]
  assign _T_5342 = ramWreqd1_6_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1585.4]
  assign _T_5346 = ramWreqd1_6_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1587.4]
  assign _T_5351 = ramWreqd1_6_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1591.4]
  assign _T_5355 = ramWreqd1_6_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1593.4]
  assign _T_5360 = ramWreqd1_6_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1597.4]
  assign _T_5364 = ramWreqd1_6_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1599.4]
  assign _T_5369 = ramWreqd1_6_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1603.4]
  assign _T_5373 = ramWreqd1_6_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1605.4]
  assign _T_5378 = ramWreqd1_7_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1609.4]
  assign _T_5382 = ramWreqd1_7_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1611.4]
  assign _T_5387 = ramWreqd1_7_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1615.4]
  assign _T_5391 = ramWreqd1_7_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1617.4]
  assign _T_5396 = ramWreqd1_7_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1621.4]
  assign _T_5400 = ramWreqd1_7_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1623.4]
  assign _T_5405 = ramWreqd1_7_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1627.4]
  assign _T_5409 = ramWreqd1_7_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1629.4]
  assign _T_5414 = ramWreqd1_8_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1633.4]
  assign _T_5418 = ramWreqd1_8_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1635.4]
  assign _T_5423 = ramWreqd1_8_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1639.4]
  assign _T_5427 = ramWreqd1_8_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1641.4]
  assign _T_5432 = ramWreqd1_8_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1645.4]
  assign _T_5436 = ramWreqd1_8_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1647.4]
  assign _T_5441 = ramWreqd1_8_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1651.4]
  assign _T_5445 = ramWreqd1_8_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1653.4]
  assign _T_5450 = ramWreqd1_9_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1657.4]
  assign _T_5454 = ramWreqd1_9_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1659.4]
  assign _T_5459 = ramWreqd1_9_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1663.4]
  assign _T_5463 = ramWreqd1_9_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1665.4]
  assign _T_5468 = ramWreqd1_9_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1669.4]
  assign _T_5472 = ramWreqd1_9_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1671.4]
  assign _T_5477 = ramWreqd1_9_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1675.4]
  assign _T_5481 = ramWreqd1_9_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1677.4]
  assign _T_5486 = ramWreqd1_10_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1681.4]
  assign _T_5490 = ramWreqd1_10_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1683.4]
  assign _T_5495 = ramWreqd1_10_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1687.4]
  assign _T_5499 = ramWreqd1_10_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1689.4]
  assign _T_5504 = ramWreqd1_10_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1693.4]
  assign _T_5508 = ramWreqd1_10_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1695.4]
  assign _T_5513 = ramWreqd1_10_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1699.4]
  assign _T_5517 = ramWreqd1_10_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1701.4]
  assign _T_5522 = ramWreqd1_11_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1705.4]
  assign _T_5526 = ramWreqd1_11_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1707.4]
  assign _T_5531 = ramWreqd1_11_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1711.4]
  assign _T_5535 = ramWreqd1_11_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1713.4]
  assign _T_5540 = ramWreqd1_11_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1717.4]
  assign _T_5544 = ramWreqd1_11_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1719.4]
  assign _T_5549 = ramWreqd1_11_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1723.4]
  assign _T_5553 = ramWreqd1_11_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1725.4]
  assign _T_5558 = ramWreqd1_12_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1729.4]
  assign _T_5562 = ramWreqd1_12_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1731.4]
  assign _T_5567 = ramWreqd1_12_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1735.4]
  assign _T_5571 = ramWreqd1_12_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1737.4]
  assign _T_5576 = ramWreqd1_12_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1741.4]
  assign _T_5580 = ramWreqd1_12_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1743.4]
  assign _T_5585 = ramWreqd1_12_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1747.4]
  assign _T_5589 = ramWreqd1_12_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1749.4]
  assign _T_5594 = ramWreqd1_13_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1753.4]
  assign _T_5598 = ramWreqd1_13_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1755.4]
  assign _T_5603 = ramWreqd1_13_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1759.4]
  assign _T_5607 = ramWreqd1_13_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1761.4]
  assign _T_5612 = ramWreqd1_13_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1765.4]
  assign _T_5616 = ramWreqd1_13_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1767.4]
  assign _T_5621 = ramWreqd1_13_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1771.4]
  assign _T_5625 = ramWreqd1_13_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1773.4]
  assign _T_5630 = ramWreqd1_14_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 105:31:@1777.4]
  assign _T_5634 = ramWreqd1_14_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 105:80:@1779.4]
  assign _T_5639 = ramWreqd1_14_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 106:31:@1783.4]
  assign _T_5643 = ramWreqd1_14_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 106:80:@1785.4]
  assign _T_5648 = ramWreqd1_14_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 107:31:@1789.4]
  assign _T_5652 = ramWreqd1_14_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 107:81:@1791.4]
  assign _T_5657 = ramWreqd1_14_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 108:31:@1795.4]
  assign _T_5661 = ramWreqd1_14_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 108:81:@1797.4]
  assign _T_10644 = io_sc2bufDat_addr[11:8]; // @[Cbuf.scala 129:28:@2524.4]
  assign datRreq_0_0 = 4'h0 == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_1_0 = 4'h1 == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_2_0 = 4'h2 == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_3_0 = 4'h3 == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_4_0 = 4'h4 == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_5_0 = 4'h5 == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_6_0 = 4'h6 == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_7_0 = 4'h7 == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_8_0 = 4'h8 == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_9_0 = 4'h9 == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_10_0 = 4'ha == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_11_0 = 4'hb == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_12_0 = 4'hc == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_13_0 = 4'hd == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign datRreq_14_0 = 4'he == _T_10644 ? io_sc2bufDat_enable : 1'h0; // @[Cbuf.scala 129:36:@2528.4]
  assign _T_10687 = io_sc2bufWt_addr[11:8]; // @[Cbuf.scala 132:26:@2535.4]
  assign wtRreq_1_0 = 4'h1 == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_2_0 = 4'h2 == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_3_0 = 4'h3 == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_4_0 = 4'h4 == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_5_0 = 4'h5 == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_6_0 = 4'h6 == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_7_0 = 4'h7 == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_8_0 = 4'h8 == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_9_0 = 4'h9 == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_10_0 = 4'ha == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_11_0 = 4'hb == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_12_0 = 4'hc == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_13_0 = 4'hd == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_14_0 = 4'he == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign wtRreq_15_0 = 4'hf == _T_10687 ? io_sc2bufWt_enable : 1'h0; // @[Cbuf.scala 132:34:@2539.4]
  assign _T_15704 = datRreq_1_0 | wtRreq_1_0; // @[Cbuf.scala 149:38:@2712.4]
  assign _T_15706 = datRreq_2_0 | wtRreq_2_0; // @[Cbuf.scala 149:38:@2716.4]
  assign _T_15708 = datRreq_3_0 | wtRreq_3_0; // @[Cbuf.scala 149:38:@2720.4]
  assign _T_15710 = datRreq_4_0 | wtRreq_4_0; // @[Cbuf.scala 149:38:@2724.4]
  assign _T_15712 = datRreq_5_0 | wtRreq_5_0; // @[Cbuf.scala 149:38:@2728.4]
  assign _T_15714 = datRreq_6_0 | wtRreq_6_0; // @[Cbuf.scala 149:38:@2732.4]
  assign _T_15716 = datRreq_7_0 | wtRreq_7_0; // @[Cbuf.scala 149:38:@2736.4]
  assign _T_15718 = datRreq_8_0 | wtRreq_8_0; // @[Cbuf.scala 149:38:@2740.4]
  assign _T_15720 = datRreq_9_0 | wtRreq_9_0; // @[Cbuf.scala 149:38:@2744.4]
  assign _T_15722 = datRreq_10_0 | wtRreq_10_0; // @[Cbuf.scala 149:38:@2748.4]
  assign _T_15724 = datRreq_11_0 | wtRreq_11_0; // @[Cbuf.scala 149:38:@2752.4]
  assign _T_15726 = datRreq_12_0 | wtRreq_12_0; // @[Cbuf.scala 149:38:@2756.4]
  assign _T_15728 = datRreq_13_0 | wtRreq_13_0; // @[Cbuf.scala 149:38:@2760.4]
  assign _T_15730 = datRreq_14_0 | wtRreq_14_0; // @[Cbuf.scala 149:38:@2764.4]
  assign _T_15732 = wtRreq_15_0 | io_sc2bufWMB_enable; // @[Cbuf.scala 145:37:@2768.4]
  assign _T_15737 = datRreq_0_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 156:28:@2773.4]
  assign _T_15745 = datRreq_1_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2779.4]
  assign _T_15749 = wtRreq_1_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2781.4]
  assign _T_15750 = _T_15745 | _T_15749; // @[Cbuf.scala 164:76:@2782.4]
  assign _T_15763 = datRreq_2_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2791.4]
  assign _T_15767 = wtRreq_2_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2793.4]
  assign _T_15768 = _T_15763 | _T_15767; // @[Cbuf.scala 164:76:@2794.4]
  assign _T_15781 = datRreq_3_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2803.4]
  assign _T_15785 = wtRreq_3_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2805.4]
  assign _T_15786 = _T_15781 | _T_15785; // @[Cbuf.scala 164:76:@2806.4]
  assign _T_15799 = datRreq_4_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2815.4]
  assign _T_15803 = wtRreq_4_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2817.4]
  assign _T_15804 = _T_15799 | _T_15803; // @[Cbuf.scala 164:76:@2818.4]
  assign _T_15817 = datRreq_5_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2827.4]
  assign _T_15821 = wtRreq_5_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2829.4]
  assign _T_15822 = _T_15817 | _T_15821; // @[Cbuf.scala 164:76:@2830.4]
  assign _T_15835 = datRreq_6_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2839.4]
  assign _T_15839 = wtRreq_6_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2841.4]
  assign _T_15840 = _T_15835 | _T_15839; // @[Cbuf.scala 164:76:@2842.4]
  assign _T_15853 = datRreq_7_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2851.4]
  assign _T_15857 = wtRreq_7_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2853.4]
  assign _T_15858 = _T_15853 | _T_15857; // @[Cbuf.scala 164:76:@2854.4]
  assign _T_15871 = datRreq_8_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2863.4]
  assign _T_15875 = wtRreq_8_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2865.4]
  assign _T_15876 = _T_15871 | _T_15875; // @[Cbuf.scala 164:76:@2866.4]
  assign _T_15889 = datRreq_9_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2875.4]
  assign _T_15893 = wtRreq_9_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2877.4]
  assign _T_15894 = _T_15889 | _T_15893; // @[Cbuf.scala 164:76:@2878.4]
  assign _T_15907 = datRreq_10_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2887.4]
  assign _T_15911 = wtRreq_10_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2889.4]
  assign _T_15912 = _T_15907 | _T_15911; // @[Cbuf.scala 164:76:@2890.4]
  assign _T_15925 = datRreq_11_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2899.4]
  assign _T_15929 = wtRreq_11_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2901.4]
  assign _T_15930 = _T_15925 | _T_15929; // @[Cbuf.scala 164:76:@2902.4]
  assign _T_15943 = datRreq_12_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2911.4]
  assign _T_15947 = wtRreq_12_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2913.4]
  assign _T_15948 = _T_15943 | _T_15947; // @[Cbuf.scala 164:76:@2914.4]
  assign _T_15961 = datRreq_13_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2923.4]
  assign _T_15965 = wtRreq_13_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2925.4]
  assign _T_15966 = _T_15961 | _T_15965; // @[Cbuf.scala 164:76:@2926.4]
  assign _T_15979 = datRreq_14_0 ? io_sc2bufDat_addr : 12'h0; // @[Cbuf.scala 164:28:@2935.4]
  assign _T_15983 = wtRreq_14_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 164:81:@2937.4]
  assign _T_15984 = _T_15979 | _T_15983; // @[Cbuf.scala 164:76:@2938.4]
  assign _T_15997 = wtRreq_15_0 ? io_sc2bufWt_addr : 12'h0; // @[Cbuf.scala 160:28:@2947.4]
  assign _T_16001 = io_sc2bufWMB_enable ? io_sc2bufWMB_addr : 12'h0; // @[Cbuf.scala 160:79:@2949.4]
  assign _T_16002 = _T_15997 | _T_16001; // @[Cbuf.scala 160:74:@2950.4]
  assign _T_26912 = datRreqd2_0_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3220.4]
  assign _T_26916 = datRreqd2_0_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3222.4]
  assign _T_26917 = {_T_26912,_T_26916}; // @[Cat.scala 30:58:@3223.4]
  assign ramdout_0_1 = RamSync_1_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3158.4 Cbuf.scala 207:21:@3563.4]
  assign ramdout_0_0 = RamSync_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3157.4 Cbuf.scala 207:21:@3556.4]
  assign _T_26918 = {ramdout_0_1,ramdout_0_0}; // @[Cat.scala 30:58:@3224.4]
  assign _T_26919 = _T_26917 & _T_26918; // @[Cbuf.scala 186:105:@3225.4]
  assign _T_26923 = datRreqd2_1_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3227.4]
  assign _T_26927 = datRreqd2_1_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3229.4]
  assign _T_26928 = {_T_26923,_T_26927}; // @[Cat.scala 30:58:@3230.4]
  assign ramdout_1_1 = RamSync_3_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3160.4 Cbuf.scala 207:21:@3577.4]
  assign ramdout_1_0 = RamSync_2_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3159.4 Cbuf.scala 207:21:@3570.4]
  assign _T_26929 = {ramdout_1_1,ramdout_1_0}; // @[Cat.scala 30:58:@3231.4]
  assign _T_26930 = _T_26928 & _T_26929; // @[Cbuf.scala 186:105:@3232.4]
  assign _T_26934 = datRreqd2_2_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3234.4]
  assign _T_26938 = datRreqd2_2_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3236.4]
  assign _T_26939 = {_T_26934,_T_26938}; // @[Cat.scala 30:58:@3237.4]
  assign ramdout_2_1 = RamSync_5_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3162.4 Cbuf.scala 207:21:@3591.4]
  assign ramdout_2_0 = RamSync_4_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3161.4 Cbuf.scala 207:21:@3584.4]
  assign _T_26940 = {ramdout_2_1,ramdout_2_0}; // @[Cat.scala 30:58:@3238.4]
  assign _T_26941 = _T_26939 & _T_26940; // @[Cbuf.scala 186:105:@3239.4]
  assign _T_26945 = datRreqd2_3_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3241.4]
  assign _T_26949 = datRreqd2_3_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3243.4]
  assign _T_26950 = {_T_26945,_T_26949}; // @[Cat.scala 30:58:@3244.4]
  assign ramdout_3_1 = RamSync_7_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3164.4 Cbuf.scala 207:21:@3605.4]
  assign ramdout_3_0 = RamSync_6_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3163.4 Cbuf.scala 207:21:@3598.4]
  assign _T_26951 = {ramdout_3_1,ramdout_3_0}; // @[Cat.scala 30:58:@3245.4]
  assign _T_26952 = _T_26950 & _T_26951; // @[Cbuf.scala 186:105:@3246.4]
  assign _T_26956 = datRreqd2_4_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3248.4]
  assign _T_26960 = datRreqd2_4_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3250.4]
  assign _T_26961 = {_T_26956,_T_26960}; // @[Cat.scala 30:58:@3251.4]
  assign ramdout_4_1 = RamSync_9_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3166.4 Cbuf.scala 207:21:@3619.4]
  assign ramdout_4_0 = RamSync_8_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3165.4 Cbuf.scala 207:21:@3612.4]
  assign _T_26962 = {ramdout_4_1,ramdout_4_0}; // @[Cat.scala 30:58:@3252.4]
  assign _T_26963 = _T_26961 & _T_26962; // @[Cbuf.scala 186:105:@3253.4]
  assign _T_26967 = datRreqd2_5_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3255.4]
  assign _T_26971 = datRreqd2_5_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3257.4]
  assign _T_26972 = {_T_26967,_T_26971}; // @[Cat.scala 30:58:@3258.4]
  assign ramdout_5_1 = RamSync_11_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3168.4 Cbuf.scala 207:21:@3633.4]
  assign ramdout_5_0 = RamSync_10_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3167.4 Cbuf.scala 207:21:@3626.4]
  assign _T_26973 = {ramdout_5_1,ramdout_5_0}; // @[Cat.scala 30:58:@3259.4]
  assign _T_26974 = _T_26972 & _T_26973; // @[Cbuf.scala 186:105:@3260.4]
  assign _T_26978 = datRreqd2_6_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3262.4]
  assign _T_26982 = datRreqd2_6_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3264.4]
  assign _T_26983 = {_T_26978,_T_26982}; // @[Cat.scala 30:58:@3265.4]
  assign ramdout_6_1 = RamSync_13_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3170.4 Cbuf.scala 207:21:@3647.4]
  assign ramdout_6_0 = RamSync_12_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3169.4 Cbuf.scala 207:21:@3640.4]
  assign _T_26984 = {ramdout_6_1,ramdout_6_0}; // @[Cat.scala 30:58:@3266.4]
  assign _T_26985 = _T_26983 & _T_26984; // @[Cbuf.scala 186:105:@3267.4]
  assign _T_26989 = datRreqd2_7_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3269.4]
  assign _T_26993 = datRreqd2_7_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3271.4]
  assign _T_26994 = {_T_26989,_T_26993}; // @[Cat.scala 30:58:@3272.4]
  assign ramdout_7_1 = RamSync_15_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3172.4 Cbuf.scala 207:21:@3661.4]
  assign ramdout_7_0 = RamSync_14_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3171.4 Cbuf.scala 207:21:@3654.4]
  assign _T_26995 = {ramdout_7_1,ramdout_7_0}; // @[Cat.scala 30:58:@3273.4]
  assign _T_26996 = _T_26994 & _T_26995; // @[Cbuf.scala 186:105:@3274.4]
  assign _T_27000 = datRreqd2_8_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3276.4]
  assign _T_27004 = datRreqd2_8_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3278.4]
  assign _T_27005 = {_T_27000,_T_27004}; // @[Cat.scala 30:58:@3279.4]
  assign ramdout_8_1 = RamSync_17_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3174.4 Cbuf.scala 207:21:@3675.4]
  assign ramdout_8_0 = RamSync_16_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3173.4 Cbuf.scala 207:21:@3668.4]
  assign _T_27006 = {ramdout_8_1,ramdout_8_0}; // @[Cat.scala 30:58:@3280.4]
  assign _T_27007 = _T_27005 & _T_27006; // @[Cbuf.scala 186:105:@3281.4]
  assign _T_27011 = datRreqd2_9_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3283.4]
  assign _T_27015 = datRreqd2_9_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3285.4]
  assign _T_27016 = {_T_27011,_T_27015}; // @[Cat.scala 30:58:@3286.4]
  assign ramdout_9_1 = RamSync_19_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3176.4 Cbuf.scala 207:21:@3689.4]
  assign ramdout_9_0 = RamSync_18_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3175.4 Cbuf.scala 207:21:@3682.4]
  assign _T_27017 = {ramdout_9_1,ramdout_9_0}; // @[Cat.scala 30:58:@3287.4]
  assign _T_27018 = _T_27016 & _T_27017; // @[Cbuf.scala 186:105:@3288.4]
  assign _T_27022 = datRreqd2_10_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3290.4]
  assign _T_27026 = datRreqd2_10_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3292.4]
  assign _T_27027 = {_T_27022,_T_27026}; // @[Cat.scala 30:58:@3293.4]
  assign ramdout_10_1 = RamSync_21_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3178.4 Cbuf.scala 207:21:@3703.4]
  assign ramdout_10_0 = RamSync_20_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3177.4 Cbuf.scala 207:21:@3696.4]
  assign _T_27028 = {ramdout_10_1,ramdout_10_0}; // @[Cat.scala 30:58:@3294.4]
  assign _T_27029 = _T_27027 & _T_27028; // @[Cbuf.scala 186:105:@3295.4]
  assign _T_27033 = datRreqd2_11_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3297.4]
  assign _T_27037 = datRreqd2_11_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3299.4]
  assign _T_27038 = {_T_27033,_T_27037}; // @[Cat.scala 30:58:@3300.4]
  assign ramdout_11_1 = RamSync_23_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3180.4 Cbuf.scala 207:21:@3717.4]
  assign ramdout_11_0 = RamSync_22_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3179.4 Cbuf.scala 207:21:@3710.4]
  assign _T_27039 = {ramdout_11_1,ramdout_11_0}; // @[Cat.scala 30:58:@3301.4]
  assign _T_27040 = _T_27038 & _T_27039; // @[Cbuf.scala 186:105:@3302.4]
  assign _T_27044 = datRreqd2_12_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3304.4]
  assign _T_27048 = datRreqd2_12_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3306.4]
  assign _T_27049 = {_T_27044,_T_27048}; // @[Cat.scala 30:58:@3307.4]
  assign ramdout_12_1 = RamSync_25_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3182.4 Cbuf.scala 207:21:@3731.4]
  assign ramdout_12_0 = RamSync_24_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3181.4 Cbuf.scala 207:21:@3724.4]
  assign _T_27050 = {ramdout_12_1,ramdout_12_0}; // @[Cat.scala 30:58:@3308.4]
  assign _T_27051 = _T_27049 & _T_27050; // @[Cbuf.scala 186:105:@3309.4]
  assign _T_27055 = datRreqd2_13_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3311.4]
  assign _T_27059 = datRreqd2_13_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3313.4]
  assign _T_27060 = {_T_27055,_T_27059}; // @[Cat.scala 30:58:@3314.4]
  assign ramdout_13_1 = RamSync_27_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3184.4 Cbuf.scala 207:21:@3745.4]
  assign ramdout_13_0 = RamSync_26_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3183.4 Cbuf.scala 207:21:@3738.4]
  assign _T_27061 = {ramdout_13_1,ramdout_13_0}; // @[Cat.scala 30:58:@3315.4]
  assign _T_27062 = _T_27060 & _T_27061; // @[Cbuf.scala 186:105:@3316.4]
  assign _T_27066 = datRreqd2_14_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3318.4]
  assign _T_27070 = datRreqd2_14_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3320.4]
  assign _T_27071 = {_T_27066,_T_27070}; // @[Cat.scala 30:58:@3321.4]
  assign ramdout_14_1 = RamSync_29_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3186.4 Cbuf.scala 207:21:@3759.4]
  assign ramdout_14_0 = RamSync_28_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3185.4 Cbuf.scala 207:21:@3752.4]
  assign _T_27072 = {ramdout_14_1,ramdout_14_0}; // @[Cat.scala 30:58:@3322.4]
  assign _T_27073 = _T_27071 & _T_27072; // @[Cbuf.scala 186:105:@3323.4]
  assign _T_27074 = _T_26919 | _T_26930; // @[Cbuf.scala 186:151:@3324.4]
  assign _T_27075 = _T_27074 | _T_26941; // @[Cbuf.scala 186:151:@3325.4]
  assign _T_27076 = _T_27075 | _T_26952; // @[Cbuf.scala 186:151:@3326.4]
  assign _T_27077 = _T_27076 | _T_26963; // @[Cbuf.scala 186:151:@3327.4]
  assign _T_27078 = _T_27077 | _T_26974; // @[Cbuf.scala 186:151:@3328.4]
  assign _T_27079 = _T_27078 | _T_26985; // @[Cbuf.scala 186:151:@3329.4]
  assign _T_27080 = _T_27079 | _T_26996; // @[Cbuf.scala 186:151:@3330.4]
  assign _T_27081 = _T_27080 | _T_27007; // @[Cbuf.scala 186:151:@3331.4]
  assign _T_27082 = _T_27081 | _T_27018; // @[Cbuf.scala 186:151:@3332.4]
  assign _T_27083 = _T_27082 | _T_27029; // @[Cbuf.scala 186:151:@3333.4]
  assign _T_27084 = _T_27083 | _T_27040; // @[Cbuf.scala 186:151:@3334.4]
  assign _T_27085 = _T_27084 | _T_27051; // @[Cbuf.scala 186:151:@3335.4]
  assign _T_27086 = _T_27085 | _T_27062; // @[Cbuf.scala 186:151:@3336.4]
  assign _T_27095 = wtRreqd2_1_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3345.4]
  assign _T_27099 = wtRreqd2_1_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3347.4]
  assign _T_27100 = {_T_27095,_T_27099}; // @[Cat.scala 30:58:@3348.4]
  assign _T_27102 = _T_27100 & _T_26929; // @[Cbuf.scala 188:103:@3350.4]
  assign _T_27106 = wtRreqd2_2_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3352.4]
  assign _T_27110 = wtRreqd2_2_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3354.4]
  assign _T_27111 = {_T_27106,_T_27110}; // @[Cat.scala 30:58:@3355.4]
  assign _T_27113 = _T_27111 & _T_26940; // @[Cbuf.scala 188:103:@3357.4]
  assign _T_27117 = wtRreqd2_3_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3359.4]
  assign _T_27121 = wtRreqd2_3_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3361.4]
  assign _T_27122 = {_T_27117,_T_27121}; // @[Cat.scala 30:58:@3362.4]
  assign _T_27124 = _T_27122 & _T_26951; // @[Cbuf.scala 188:103:@3364.4]
  assign _T_27128 = wtRreqd2_4_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3366.4]
  assign _T_27132 = wtRreqd2_4_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3368.4]
  assign _T_27133 = {_T_27128,_T_27132}; // @[Cat.scala 30:58:@3369.4]
  assign _T_27135 = _T_27133 & _T_26962; // @[Cbuf.scala 188:103:@3371.4]
  assign _T_27139 = wtRreqd2_5_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3373.4]
  assign _T_27143 = wtRreqd2_5_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3375.4]
  assign _T_27144 = {_T_27139,_T_27143}; // @[Cat.scala 30:58:@3376.4]
  assign _T_27146 = _T_27144 & _T_26973; // @[Cbuf.scala 188:103:@3378.4]
  assign _T_27150 = wtRreqd2_6_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3380.4]
  assign _T_27154 = wtRreqd2_6_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3382.4]
  assign _T_27155 = {_T_27150,_T_27154}; // @[Cat.scala 30:58:@3383.4]
  assign _T_27157 = _T_27155 & _T_26984; // @[Cbuf.scala 188:103:@3385.4]
  assign _T_27161 = wtRreqd2_7_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3387.4]
  assign _T_27165 = wtRreqd2_7_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3389.4]
  assign _T_27166 = {_T_27161,_T_27165}; // @[Cat.scala 30:58:@3390.4]
  assign _T_27168 = _T_27166 & _T_26995; // @[Cbuf.scala 188:103:@3392.4]
  assign _T_27172 = wtRreqd2_8_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3394.4]
  assign _T_27176 = wtRreqd2_8_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3396.4]
  assign _T_27177 = {_T_27172,_T_27176}; // @[Cat.scala 30:58:@3397.4]
  assign _T_27179 = _T_27177 & _T_27006; // @[Cbuf.scala 188:103:@3399.4]
  assign _T_27183 = wtRreqd2_9_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3401.4]
  assign _T_27187 = wtRreqd2_9_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3403.4]
  assign _T_27188 = {_T_27183,_T_27187}; // @[Cat.scala 30:58:@3404.4]
  assign _T_27190 = _T_27188 & _T_27017; // @[Cbuf.scala 188:103:@3406.4]
  assign _T_27194 = wtRreqd2_10_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3408.4]
  assign _T_27198 = wtRreqd2_10_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3410.4]
  assign _T_27199 = {_T_27194,_T_27198}; // @[Cat.scala 30:58:@3411.4]
  assign _T_27201 = _T_27199 & _T_27028; // @[Cbuf.scala 188:103:@3413.4]
  assign _T_27205 = wtRreqd2_11_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3415.4]
  assign _T_27209 = wtRreqd2_11_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3417.4]
  assign _T_27210 = {_T_27205,_T_27209}; // @[Cat.scala 30:58:@3418.4]
  assign _T_27212 = _T_27210 & _T_27039; // @[Cbuf.scala 188:103:@3420.4]
  assign _T_27216 = wtRreqd2_12_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3422.4]
  assign _T_27220 = wtRreqd2_12_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3424.4]
  assign _T_27221 = {_T_27216,_T_27220}; // @[Cat.scala 30:58:@3425.4]
  assign _T_27223 = _T_27221 & _T_27050; // @[Cbuf.scala 188:103:@3427.4]
  assign _T_27227 = wtRreqd2_13_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3429.4]
  assign _T_27231 = wtRreqd2_13_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3431.4]
  assign _T_27232 = {_T_27227,_T_27231}; // @[Cat.scala 30:58:@3432.4]
  assign _T_27234 = _T_27232 & _T_27061; // @[Cbuf.scala 188:103:@3434.4]
  assign _T_27238 = wtRreqd2_14_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3436.4]
  assign _T_27242 = wtRreqd2_14_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3438.4]
  assign _T_27243 = {_T_27238,_T_27242}; // @[Cat.scala 30:58:@3439.4]
  assign _T_27245 = _T_27243 & _T_27072; // @[Cbuf.scala 188:103:@3441.4]
  assign _T_27249 = wtRreqd2_15_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3443.4]
  assign _T_27253 = wtRreqd2_15_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3445.4]
  assign _T_27254 = {_T_27249,_T_27253}; // @[Cat.scala 30:58:@3446.4]
  assign ramdout_15_1 = RamSync_31_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3188.4 Cbuf.scala 207:21:@3773.4]
  assign ramdout_15_0 = RamSync_30_io_dout; // @[Cbuf.scala 174:24:@3156.4 Cbuf.scala 174:24:@3187.4 Cbuf.scala 207:21:@3766.4]
  assign _T_27255 = {ramdout_15_1,ramdout_15_0}; // @[Cat.scala 30:58:@3447.4]
  assign _T_27256 = _T_27254 & _T_27255; // @[Cbuf.scala 188:103:@3448.4]
  assign _T_27257 = _T_27102 | _T_27113; // @[Cbuf.scala 188:149:@3449.4]
  assign _T_27258 = _T_27257 | _T_27124; // @[Cbuf.scala 188:149:@3450.4]
  assign _T_27259 = _T_27258 | _T_27135; // @[Cbuf.scala 188:149:@3451.4]
  assign _T_27260 = _T_27259 | _T_27146; // @[Cbuf.scala 188:149:@3452.4]
  assign _T_27261 = _T_27260 | _T_27157; // @[Cbuf.scala 188:149:@3453.4]
  assign _T_27262 = _T_27261 | _T_27168; // @[Cbuf.scala 188:149:@3454.4]
  assign _T_27263 = _T_27262 | _T_27179; // @[Cbuf.scala 188:149:@3455.4]
  assign _T_27264 = _T_27263 | _T_27190; // @[Cbuf.scala 188:149:@3456.4]
  assign _T_27265 = _T_27264 | _T_27201; // @[Cbuf.scala 188:149:@3457.4]
  assign _T_27266 = _T_27265 | _T_27212; // @[Cbuf.scala 188:149:@3458.4]
  assign _T_27267 = _T_27266 | _T_27223; // @[Cbuf.scala 188:149:@3459.4]
  assign _T_27268 = _T_27267 | _T_27234; // @[Cbuf.scala 188:149:@3460.4]
  assign _T_27269 = _T_27268 | _T_27245; // @[Cbuf.scala 188:149:@3461.4]
  assign _T_27278 = wmbRreqd2_1 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3470.4]
  assign _T_27282 = wmbRreqd2_0 ? 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 512'h0; // @[Bitwise.scala 72:12:@3472.4]
  assign _T_27283 = {_T_27278,_T_27282}; // @[Cat.scala 30:58:@3473.4]
  assign io_sc2bufDat_data = p0Datad6; // @[Cbuf.scala 216:21:@3778.4]
  assign io_sc2bufDat_valid = p0Validd6; // @[Cbuf.scala 217:22:@3779.4]
  assign io_sc2bufWt_data = p1Datad6; // @[Cbuf.scala 218:20:@3780.4]
  assign io_sc2bufWt_valid = p1Validd6; // @[Cbuf.scala 219:21:@3781.4]
  assign io_sc2bufWMB_data = p2Datad6; // @[Cbuf.scala 220:21:@3782.4]
  assign io_sc2bufWMB_valid = p2Validd6; // @[Cbuf.scala 221:22:@3783.4]
  assign RamSync_clock = clock; // @[:@649.4]
  assign RamSync_io_re = ramRreq_0_0; // @[Cbuf.scala 205:24:@3554.4]
  assign RamSync_io_we = ramWreqd2_0_0; // @[Cbuf.scala 209:24:@3557.4]
  assign RamSync_io_ra = ramRaddr_0_0; // @[Cbuf.scala 206:24:@3555.4]
  assign RamSync_io_wa = ramWreqd1_0_0 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 210:24:@3558.4]
  assign RamSync_io_di = ramWreqd1_0_0 ? ramp0DatLod1 : 512'h0; // @[Cbuf.scala 211:24:@3559.4]
  assign RamSync_1_clock = clock; // @[:@652.4]
  assign RamSync_1_io_re = ramRreq_0_1; // @[Cbuf.scala 205:24:@3561.4]
  assign RamSync_1_io_we = ramWreqd2_0_1; // @[Cbuf.scala 209:24:@3564.4]
  assign RamSync_1_io_ra = ramRaddr_0_1; // @[Cbuf.scala 206:24:@3562.4]
  assign RamSync_1_io_wa = ramWreqd1_0_1 ? ramp0Addrd1 : 8'h0; // @[Cbuf.scala 210:24:@3565.4]
  assign RamSync_1_io_di = ramWreqd1_0_1 ? ramp0DatHid1 : 512'h0; // @[Cbuf.scala 211:24:@3566.4]
  assign RamSync_2_clock = clock; // @[:@655.4]
  assign RamSync_2_io_re = ramRreq_1_0; // @[Cbuf.scala 205:24:@3568.4]
  assign RamSync_2_io_we = ramWreqd2_1_0; // @[Cbuf.scala 209:24:@3571.4]
  assign RamSync_2_io_ra = ramRaddr_1_0; // @[Cbuf.scala 206:24:@3569.4]
  assign RamSync_2_io_wa = _T_5162 | _T_5166; // @[Cbuf.scala 210:24:@3572.4]
  assign RamSync_2_io_di = _T_5180 | _T_5184; // @[Cbuf.scala 211:24:@3573.4]
  assign RamSync_3_clock = clock; // @[:@658.4]
  assign RamSync_3_io_re = ramRreq_1_1; // @[Cbuf.scala 205:24:@3575.4]
  assign RamSync_3_io_we = ramWreqd2_1_1; // @[Cbuf.scala 209:24:@3578.4]
  assign RamSync_3_io_ra = ramRaddr_1_1; // @[Cbuf.scala 206:24:@3576.4]
  assign RamSync_3_io_wa = _T_5171 | _T_5175; // @[Cbuf.scala 210:24:@3579.4]
  assign RamSync_3_io_di = _T_5189 | _T_5193; // @[Cbuf.scala 211:24:@3580.4]
  assign RamSync_4_clock = clock; // @[:@661.4]
  assign RamSync_4_io_re = ramRreq_2_0; // @[Cbuf.scala 205:24:@3582.4]
  assign RamSync_4_io_we = ramWreqd2_2_0; // @[Cbuf.scala 209:24:@3585.4]
  assign RamSync_4_io_ra = ramRaddr_2_0; // @[Cbuf.scala 206:24:@3583.4]
  assign RamSync_4_io_wa = _T_5198 | _T_5202; // @[Cbuf.scala 210:24:@3586.4]
  assign RamSync_4_io_di = _T_5216 | _T_5220; // @[Cbuf.scala 211:24:@3587.4]
  assign RamSync_5_clock = clock; // @[:@664.4]
  assign RamSync_5_io_re = ramRreq_2_1; // @[Cbuf.scala 205:24:@3589.4]
  assign RamSync_5_io_we = ramWreqd2_2_1; // @[Cbuf.scala 209:24:@3592.4]
  assign RamSync_5_io_ra = ramRaddr_2_1; // @[Cbuf.scala 206:24:@3590.4]
  assign RamSync_5_io_wa = _T_5207 | _T_5211; // @[Cbuf.scala 210:24:@3593.4]
  assign RamSync_5_io_di = _T_5225 | _T_5229; // @[Cbuf.scala 211:24:@3594.4]
  assign RamSync_6_clock = clock; // @[:@667.4]
  assign RamSync_6_io_re = ramRreq_3_0; // @[Cbuf.scala 205:24:@3596.4]
  assign RamSync_6_io_we = ramWreqd2_3_0; // @[Cbuf.scala 209:24:@3599.4]
  assign RamSync_6_io_ra = ramRaddr_3_0; // @[Cbuf.scala 206:24:@3597.4]
  assign RamSync_6_io_wa = _T_5234 | _T_5238; // @[Cbuf.scala 210:24:@3600.4]
  assign RamSync_6_io_di = _T_5252 | _T_5256; // @[Cbuf.scala 211:24:@3601.4]
  assign RamSync_7_clock = clock; // @[:@670.4]
  assign RamSync_7_io_re = ramRreq_3_1; // @[Cbuf.scala 205:24:@3603.4]
  assign RamSync_7_io_we = ramWreqd2_3_1; // @[Cbuf.scala 209:24:@3606.4]
  assign RamSync_7_io_ra = ramRaddr_3_1; // @[Cbuf.scala 206:24:@3604.4]
  assign RamSync_7_io_wa = _T_5243 | _T_5247; // @[Cbuf.scala 210:24:@3607.4]
  assign RamSync_7_io_di = _T_5261 | _T_5265; // @[Cbuf.scala 211:24:@3608.4]
  assign RamSync_8_clock = clock; // @[:@673.4]
  assign RamSync_8_io_re = ramRreq_4_0; // @[Cbuf.scala 205:24:@3610.4]
  assign RamSync_8_io_we = ramWreqd2_4_0; // @[Cbuf.scala 209:24:@3613.4]
  assign RamSync_8_io_ra = ramRaddr_4_0; // @[Cbuf.scala 206:24:@3611.4]
  assign RamSync_8_io_wa = _T_5270 | _T_5274; // @[Cbuf.scala 210:24:@3614.4]
  assign RamSync_8_io_di = _T_5288 | _T_5292; // @[Cbuf.scala 211:24:@3615.4]
  assign RamSync_9_clock = clock; // @[:@676.4]
  assign RamSync_9_io_re = ramRreq_4_1; // @[Cbuf.scala 205:24:@3617.4]
  assign RamSync_9_io_we = ramWreqd2_4_1; // @[Cbuf.scala 209:24:@3620.4]
  assign RamSync_9_io_ra = ramRaddr_4_1; // @[Cbuf.scala 206:24:@3618.4]
  assign RamSync_9_io_wa = _T_5279 | _T_5283; // @[Cbuf.scala 210:24:@3621.4]
  assign RamSync_9_io_di = _T_5297 | _T_5301; // @[Cbuf.scala 211:24:@3622.4]
  assign RamSync_10_clock = clock; // @[:@679.4]
  assign RamSync_10_io_re = ramRreq_5_0; // @[Cbuf.scala 205:24:@3624.4]
  assign RamSync_10_io_we = ramWreqd2_5_0; // @[Cbuf.scala 209:24:@3627.4]
  assign RamSync_10_io_ra = ramRaddr_5_0; // @[Cbuf.scala 206:24:@3625.4]
  assign RamSync_10_io_wa = _T_5306 | _T_5310; // @[Cbuf.scala 210:24:@3628.4]
  assign RamSync_10_io_di = _T_5324 | _T_5328; // @[Cbuf.scala 211:24:@3629.4]
  assign RamSync_11_clock = clock; // @[:@682.4]
  assign RamSync_11_io_re = ramRreq_5_1; // @[Cbuf.scala 205:24:@3631.4]
  assign RamSync_11_io_we = ramWreqd2_5_1; // @[Cbuf.scala 209:24:@3634.4]
  assign RamSync_11_io_ra = ramRaddr_5_1; // @[Cbuf.scala 206:24:@3632.4]
  assign RamSync_11_io_wa = _T_5315 | _T_5319; // @[Cbuf.scala 210:24:@3635.4]
  assign RamSync_11_io_di = _T_5333 | _T_5337; // @[Cbuf.scala 211:24:@3636.4]
  assign RamSync_12_clock = clock; // @[:@685.4]
  assign RamSync_12_io_re = ramRreq_6_0; // @[Cbuf.scala 205:24:@3638.4]
  assign RamSync_12_io_we = ramWreqd2_6_0; // @[Cbuf.scala 209:24:@3641.4]
  assign RamSync_12_io_ra = ramRaddr_6_0; // @[Cbuf.scala 206:24:@3639.4]
  assign RamSync_12_io_wa = _T_5342 | _T_5346; // @[Cbuf.scala 210:24:@3642.4]
  assign RamSync_12_io_di = _T_5360 | _T_5364; // @[Cbuf.scala 211:24:@3643.4]
  assign RamSync_13_clock = clock; // @[:@688.4]
  assign RamSync_13_io_re = ramRreq_6_1; // @[Cbuf.scala 205:24:@3645.4]
  assign RamSync_13_io_we = ramWreqd2_6_1; // @[Cbuf.scala 209:24:@3648.4]
  assign RamSync_13_io_ra = ramRaddr_6_1; // @[Cbuf.scala 206:24:@3646.4]
  assign RamSync_13_io_wa = _T_5351 | _T_5355; // @[Cbuf.scala 210:24:@3649.4]
  assign RamSync_13_io_di = _T_5369 | _T_5373; // @[Cbuf.scala 211:24:@3650.4]
  assign RamSync_14_clock = clock; // @[:@691.4]
  assign RamSync_14_io_re = ramRreq_7_0; // @[Cbuf.scala 205:24:@3652.4]
  assign RamSync_14_io_we = ramWreqd2_7_0; // @[Cbuf.scala 209:24:@3655.4]
  assign RamSync_14_io_ra = ramRaddr_7_0; // @[Cbuf.scala 206:24:@3653.4]
  assign RamSync_14_io_wa = _T_5378 | _T_5382; // @[Cbuf.scala 210:24:@3656.4]
  assign RamSync_14_io_di = _T_5396 | _T_5400; // @[Cbuf.scala 211:24:@3657.4]
  assign RamSync_15_clock = clock; // @[:@694.4]
  assign RamSync_15_io_re = ramRreq_7_1; // @[Cbuf.scala 205:24:@3659.4]
  assign RamSync_15_io_we = ramWreqd2_7_1; // @[Cbuf.scala 209:24:@3662.4]
  assign RamSync_15_io_ra = ramRaddr_7_1; // @[Cbuf.scala 206:24:@3660.4]
  assign RamSync_15_io_wa = _T_5387 | _T_5391; // @[Cbuf.scala 210:24:@3663.4]
  assign RamSync_15_io_di = _T_5405 | _T_5409; // @[Cbuf.scala 211:24:@3664.4]
  assign RamSync_16_clock = clock; // @[:@697.4]
  assign RamSync_16_io_re = ramRreq_8_0; // @[Cbuf.scala 205:24:@3666.4]
  assign RamSync_16_io_we = ramWreqd2_8_0; // @[Cbuf.scala 209:24:@3669.4]
  assign RamSync_16_io_ra = ramRaddr_8_0; // @[Cbuf.scala 206:24:@3667.4]
  assign RamSync_16_io_wa = _T_5414 | _T_5418; // @[Cbuf.scala 210:24:@3670.4]
  assign RamSync_16_io_di = _T_5432 | _T_5436; // @[Cbuf.scala 211:24:@3671.4]
  assign RamSync_17_clock = clock; // @[:@700.4]
  assign RamSync_17_io_re = ramRreq_8_1; // @[Cbuf.scala 205:24:@3673.4]
  assign RamSync_17_io_we = ramWreqd2_8_1; // @[Cbuf.scala 209:24:@3676.4]
  assign RamSync_17_io_ra = ramRaddr_8_1; // @[Cbuf.scala 206:24:@3674.4]
  assign RamSync_17_io_wa = _T_5423 | _T_5427; // @[Cbuf.scala 210:24:@3677.4]
  assign RamSync_17_io_di = _T_5441 | _T_5445; // @[Cbuf.scala 211:24:@3678.4]
  assign RamSync_18_clock = clock; // @[:@703.4]
  assign RamSync_18_io_re = ramRreq_9_0; // @[Cbuf.scala 205:24:@3680.4]
  assign RamSync_18_io_we = ramWreqd2_9_0; // @[Cbuf.scala 209:24:@3683.4]
  assign RamSync_18_io_ra = ramRaddr_9_0; // @[Cbuf.scala 206:24:@3681.4]
  assign RamSync_18_io_wa = _T_5450 | _T_5454; // @[Cbuf.scala 210:24:@3684.4]
  assign RamSync_18_io_di = _T_5468 | _T_5472; // @[Cbuf.scala 211:24:@3685.4]
  assign RamSync_19_clock = clock; // @[:@706.4]
  assign RamSync_19_io_re = ramRreq_9_1; // @[Cbuf.scala 205:24:@3687.4]
  assign RamSync_19_io_we = ramWreqd2_9_1; // @[Cbuf.scala 209:24:@3690.4]
  assign RamSync_19_io_ra = ramRaddr_9_1; // @[Cbuf.scala 206:24:@3688.4]
  assign RamSync_19_io_wa = _T_5459 | _T_5463; // @[Cbuf.scala 210:24:@3691.4]
  assign RamSync_19_io_di = _T_5477 | _T_5481; // @[Cbuf.scala 211:24:@3692.4]
  assign RamSync_20_clock = clock; // @[:@709.4]
  assign RamSync_20_io_re = ramRreq_10_0; // @[Cbuf.scala 205:24:@3694.4]
  assign RamSync_20_io_we = ramWreqd2_10_0; // @[Cbuf.scala 209:24:@3697.4]
  assign RamSync_20_io_ra = ramRaddr_10_0; // @[Cbuf.scala 206:24:@3695.4]
  assign RamSync_20_io_wa = _T_5486 | _T_5490; // @[Cbuf.scala 210:24:@3698.4]
  assign RamSync_20_io_di = _T_5504 | _T_5508; // @[Cbuf.scala 211:24:@3699.4]
  assign RamSync_21_clock = clock; // @[:@712.4]
  assign RamSync_21_io_re = ramRreq_10_1; // @[Cbuf.scala 205:24:@3701.4]
  assign RamSync_21_io_we = ramWreqd2_10_1; // @[Cbuf.scala 209:24:@3704.4]
  assign RamSync_21_io_ra = ramRaddr_10_1; // @[Cbuf.scala 206:24:@3702.4]
  assign RamSync_21_io_wa = _T_5495 | _T_5499; // @[Cbuf.scala 210:24:@3705.4]
  assign RamSync_21_io_di = _T_5513 | _T_5517; // @[Cbuf.scala 211:24:@3706.4]
  assign RamSync_22_clock = clock; // @[:@715.4]
  assign RamSync_22_io_re = ramRreq_11_0; // @[Cbuf.scala 205:24:@3708.4]
  assign RamSync_22_io_we = ramWreqd2_11_0; // @[Cbuf.scala 209:24:@3711.4]
  assign RamSync_22_io_ra = ramRaddr_11_0; // @[Cbuf.scala 206:24:@3709.4]
  assign RamSync_22_io_wa = _T_5522 | _T_5526; // @[Cbuf.scala 210:24:@3712.4]
  assign RamSync_22_io_di = _T_5540 | _T_5544; // @[Cbuf.scala 211:24:@3713.4]
  assign RamSync_23_clock = clock; // @[:@718.4]
  assign RamSync_23_io_re = ramRreq_11_1; // @[Cbuf.scala 205:24:@3715.4]
  assign RamSync_23_io_we = ramWreqd2_11_1; // @[Cbuf.scala 209:24:@3718.4]
  assign RamSync_23_io_ra = ramRaddr_11_1; // @[Cbuf.scala 206:24:@3716.4]
  assign RamSync_23_io_wa = _T_5531 | _T_5535; // @[Cbuf.scala 210:24:@3719.4]
  assign RamSync_23_io_di = _T_5549 | _T_5553; // @[Cbuf.scala 211:24:@3720.4]
  assign RamSync_24_clock = clock; // @[:@721.4]
  assign RamSync_24_io_re = ramRreq_12_0; // @[Cbuf.scala 205:24:@3722.4]
  assign RamSync_24_io_we = ramWreqd2_12_0; // @[Cbuf.scala 209:24:@3725.4]
  assign RamSync_24_io_ra = ramRaddr_12_0; // @[Cbuf.scala 206:24:@3723.4]
  assign RamSync_24_io_wa = _T_5558 | _T_5562; // @[Cbuf.scala 210:24:@3726.4]
  assign RamSync_24_io_di = _T_5576 | _T_5580; // @[Cbuf.scala 211:24:@3727.4]
  assign RamSync_25_clock = clock; // @[:@724.4]
  assign RamSync_25_io_re = ramRreq_12_1; // @[Cbuf.scala 205:24:@3729.4]
  assign RamSync_25_io_we = ramWreqd2_12_1; // @[Cbuf.scala 209:24:@3732.4]
  assign RamSync_25_io_ra = ramRaddr_12_1; // @[Cbuf.scala 206:24:@3730.4]
  assign RamSync_25_io_wa = _T_5567 | _T_5571; // @[Cbuf.scala 210:24:@3733.4]
  assign RamSync_25_io_di = _T_5585 | _T_5589; // @[Cbuf.scala 211:24:@3734.4]
  assign RamSync_26_clock = clock; // @[:@727.4]
  assign RamSync_26_io_re = ramRreq_13_0; // @[Cbuf.scala 205:24:@3736.4]
  assign RamSync_26_io_we = ramWreqd2_13_0; // @[Cbuf.scala 209:24:@3739.4]
  assign RamSync_26_io_ra = ramRaddr_13_0; // @[Cbuf.scala 206:24:@3737.4]
  assign RamSync_26_io_wa = _T_5594 | _T_5598; // @[Cbuf.scala 210:24:@3740.4]
  assign RamSync_26_io_di = _T_5612 | _T_5616; // @[Cbuf.scala 211:24:@3741.4]
  assign RamSync_27_clock = clock; // @[:@730.4]
  assign RamSync_27_io_re = ramRreq_13_1; // @[Cbuf.scala 205:24:@3743.4]
  assign RamSync_27_io_we = ramWreqd2_13_1; // @[Cbuf.scala 209:24:@3746.4]
  assign RamSync_27_io_ra = ramRaddr_13_1; // @[Cbuf.scala 206:24:@3744.4]
  assign RamSync_27_io_wa = _T_5603 | _T_5607; // @[Cbuf.scala 210:24:@3747.4]
  assign RamSync_27_io_di = _T_5621 | _T_5625; // @[Cbuf.scala 211:24:@3748.4]
  assign RamSync_28_clock = clock; // @[:@733.4]
  assign RamSync_28_io_re = ramRreq_14_0; // @[Cbuf.scala 205:24:@3750.4]
  assign RamSync_28_io_we = ramWreqd2_14_0; // @[Cbuf.scala 209:24:@3753.4]
  assign RamSync_28_io_ra = ramRaddr_14_0; // @[Cbuf.scala 206:24:@3751.4]
  assign RamSync_28_io_wa = _T_5630 | _T_5634; // @[Cbuf.scala 210:24:@3754.4]
  assign RamSync_28_io_di = _T_5648 | _T_5652; // @[Cbuf.scala 211:24:@3755.4]
  assign RamSync_29_clock = clock; // @[:@736.4]
  assign RamSync_29_io_re = ramRreq_14_1; // @[Cbuf.scala 205:24:@3757.4]
  assign RamSync_29_io_we = ramWreqd2_14_1; // @[Cbuf.scala 209:24:@3760.4]
  assign RamSync_29_io_ra = ramRaddr_14_1; // @[Cbuf.scala 206:24:@3758.4]
  assign RamSync_29_io_wa = _T_5639 | _T_5643; // @[Cbuf.scala 210:24:@3761.4]
  assign RamSync_29_io_di = _T_5657 | _T_5661; // @[Cbuf.scala 211:24:@3762.4]
  assign RamSync_30_clock = clock; // @[:@739.4]
  assign RamSync_30_io_re = ramRreq_15_0; // @[Cbuf.scala 205:24:@3764.4]
  assign RamSync_30_io_we = ramWreqd2_15_0; // @[Cbuf.scala 209:24:@3767.4]
  assign RamSync_30_io_ra = ramRaddr_15_0; // @[Cbuf.scala 206:24:@3765.4]
  assign RamSync_30_io_wa = ramWreqd1_15_0 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 210:24:@3768.4]
  assign RamSync_30_io_di = ramWreqd1_15_0 ? ramp1WtLod1 : 512'h0; // @[Cbuf.scala 211:24:@3769.4]
  assign RamSync_31_clock = clock; // @[:@742.4]
  assign RamSync_31_io_re = ramRreq_15_1; // @[Cbuf.scala 205:24:@3771.4]
  assign RamSync_31_io_we = ramWreqd2_15_1; // @[Cbuf.scala 209:24:@3774.4]
  assign RamSync_31_io_ra = ramRaddr_15_1; // @[Cbuf.scala 206:24:@3772.4]
  assign RamSync_31_io_wa = ramWreqd1_15_1 ? ramp1Addrd1 : 8'h0; // @[Cbuf.scala 210:24:@3775.4]
  assign RamSync_31_io_di = ramWreqd1_15_1 ? ramp1WtHid1 : 512'h0; // @[Cbuf.scala 211:24:@3776.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ramWreqd1_0_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ramWreqd1_0_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ramWreqd1_1_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ramWreqd1_1_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ramWreqd1_2_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ramWreqd1_2_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ramWreqd1_3_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ramWreqd1_3_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ramWreqd1_4_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  ramWreqd1_4_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  ramWreqd1_5_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  ramWreqd1_5_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  ramWreqd1_6_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  ramWreqd1_6_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  ramWreqd1_7_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  ramWreqd1_7_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  ramWreqd1_8_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  ramWreqd1_8_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  ramWreqd1_9_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  ramWreqd1_9_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  ramWreqd1_10_0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  ramWreqd1_10_1 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  ramWreqd1_11_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  ramWreqd1_11_1 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  ramWreqd1_12_0 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  ramWreqd1_12_1 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  ramWreqd1_13_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  ramWreqd1_13_1 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  ramWreqd1_14_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  ramWreqd1_14_1 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  ramWreqd1_15_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  ramWreqd1_15_1 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  ramp0Addrd1 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  ramp1Addrd1 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {16{`RANDOM}};
  ramp0DatLod1 = _RAND_34[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {16{`RANDOM}};
  ramp0DatHid1 = _RAND_35[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {16{`RANDOM}};
  ramp1WtLod1 = _RAND_36[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {16{`RANDOM}};
  ramp1WtHid1 = _RAND_37[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  ramWreqd2_0_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  ramWreqd2_0_1 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  ramWreqd2_1_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  ramWreqd2_1_1 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  ramWreqd2_2_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  ramWreqd2_2_1 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  ramWreqd2_3_0 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  ramWreqd2_3_1 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  ramWreqd2_4_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  ramWreqd2_4_1 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  ramWreqd2_5_0 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  ramWreqd2_5_1 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  ramWreqd2_6_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  ramWreqd2_6_1 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  ramWreqd2_7_0 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  ramWreqd2_7_1 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  ramWreqd2_8_0 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  ramWreqd2_8_1 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  ramWreqd2_9_0 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  ramWreqd2_9_1 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  ramWreqd2_10_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  ramWreqd2_10_1 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  ramWreqd2_11_0 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  ramWreqd2_11_1 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  ramWreqd2_12_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  ramWreqd2_12_1 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  ramWreqd2_13_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  ramWreqd2_13_1 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  ramWreqd2_14_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  ramWreqd2_14_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  ramWreqd2_15_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  ramWreqd2_15_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  ramRreq_0_0 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  ramRreq_0_1 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  ramRreq_1_0 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  ramRreq_1_1 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  ramRreq_2_0 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  ramRreq_2_1 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  ramRreq_3_0 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  ramRreq_3_1 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  ramRreq_4_0 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  ramRreq_4_1 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  ramRreq_5_0 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  ramRreq_5_1 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  ramRreq_6_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  ramRreq_6_1 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  ramRreq_7_0 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  ramRreq_7_1 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  ramRreq_8_0 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  ramRreq_8_1 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  ramRreq_9_0 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  ramRreq_9_1 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  ramRreq_10_0 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  ramRreq_10_1 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  ramRreq_11_0 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  ramRreq_11_1 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  ramRreq_12_0 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  ramRreq_12_1 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  ramRreq_13_0 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  ramRreq_13_1 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  ramRreq_14_0 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  ramRreq_14_1 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  ramRreq_15_0 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  ramRreq_15_1 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  ramRaddr_0_0 = _RAND_102[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  ramRaddr_0_1 = _RAND_103[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  ramRaddr_1_0 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  ramRaddr_1_1 = _RAND_105[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  ramRaddr_2_0 = _RAND_106[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  ramRaddr_2_1 = _RAND_107[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  ramRaddr_3_0 = _RAND_108[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  ramRaddr_3_1 = _RAND_109[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  ramRaddr_4_0 = _RAND_110[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  ramRaddr_4_1 = _RAND_111[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  ramRaddr_5_0 = _RAND_112[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  ramRaddr_5_1 = _RAND_113[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  ramRaddr_6_0 = _RAND_114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  ramRaddr_6_1 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  ramRaddr_7_0 = _RAND_116[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  ramRaddr_7_1 = _RAND_117[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  ramRaddr_8_0 = _RAND_118[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  ramRaddr_8_1 = _RAND_119[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  ramRaddr_9_0 = _RAND_120[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  ramRaddr_9_1 = _RAND_121[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  ramRaddr_10_0 = _RAND_122[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  ramRaddr_10_1 = _RAND_123[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  ramRaddr_11_0 = _RAND_124[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  ramRaddr_11_1 = _RAND_125[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  ramRaddr_12_0 = _RAND_126[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  ramRaddr_12_1 = _RAND_127[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  ramRaddr_13_0 = _RAND_128[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  ramRaddr_13_1 = _RAND_129[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  ramRaddr_14_0 = _RAND_130[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  ramRaddr_14_1 = _RAND_131[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  ramRaddr_15_0 = _RAND_132[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  ramRaddr_15_1 = _RAND_133[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_16712_0_0 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_16712_0_1 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_16712_1_0 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_16712_1_1 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_16712_2_0 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_16712_2_1 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_16712_3_0 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_16712_3_1 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_16712_4_0 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_16712_4_1 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_16712_5_0 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_16712_5_1 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_16712_6_0 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_16712_6_1 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_16712_7_0 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_16712_7_1 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_16712_8_0 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_16712_8_1 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_16712_9_0 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_16712_9_1 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_16712_10_0 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_16712_10_1 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_16712_11_0 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_16712_11_1 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_16712_12_0 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_16712_12_1 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_16712_13_0 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_16712_13_1 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_16712_14_0 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_16712_14_1 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  datRreqd2_0_0 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  datRreqd2_0_1 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  datRreqd2_1_0 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  datRreqd2_1_1 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  datRreqd2_2_0 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  datRreqd2_2_1 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  datRreqd2_3_0 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  datRreqd2_3_1 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  datRreqd2_4_0 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  datRreqd2_4_1 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  datRreqd2_5_0 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  datRreqd2_5_1 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  datRreqd2_6_0 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  datRreqd2_6_1 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  datRreqd2_7_0 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  datRreqd2_7_1 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  datRreqd2_8_0 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  datRreqd2_8_1 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  datRreqd2_9_0 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  datRreqd2_9_1 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  datRreqd2_10_0 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  datRreqd2_10_1 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  datRreqd2_11_0 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  datRreqd2_11_1 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  datRreqd2_12_0 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  datRreqd2_12_1 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  datRreqd2_13_0 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  datRreqd2_13_1 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  datRreqd2_14_0 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  datRreqd2_14_1 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_21752_1_0 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_21752_1_1 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_21752_2_0 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_21752_2_1 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_21752_3_0 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_21752_3_1 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_21752_4_0 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_21752_4_1 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_21752_5_0 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_21752_5_1 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_21752_6_0 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_21752_6_1 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_21752_7_0 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_21752_7_1 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_21752_8_0 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_21752_8_1 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_21752_9_0 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_21752_9_1 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_21752_10_0 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_21752_10_1 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_21752_11_0 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_21752_11_1 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_21752_12_0 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_21752_12_1 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_21752_13_0 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_21752_13_1 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_21752_14_0 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_21752_14_1 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_21752_15_0 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_21752_15_1 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  wtRreqd2_1_0 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  wtRreqd2_1_1 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  wtRreqd2_2_0 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  wtRreqd2_2_1 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  wtRreqd2_3_0 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  wtRreqd2_3_1 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  wtRreqd2_4_0 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  wtRreqd2_4_1 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  wtRreqd2_5_0 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  wtRreqd2_5_1 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  wtRreqd2_6_0 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  wtRreqd2_6_1 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  wtRreqd2_7_0 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  wtRreqd2_7_1 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  wtRreqd2_8_0 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  wtRreqd2_8_1 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  wtRreqd2_9_0 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  wtRreqd2_9_1 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  wtRreqd2_10_0 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  wtRreqd2_10_1 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  wtRreqd2_11_0 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  wtRreqd2_11_1 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  wtRreqd2_12_0 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  wtRreqd2_12_1 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  wtRreqd2_13_0 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  wtRreqd2_13_1 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  wtRreqd2_14_0 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  wtRreqd2_14_1 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  wtRreqd2_15_0 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  wtRreqd2_15_1 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_26101_0 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_26101_1 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  wmbRreqd2_0 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  wmbRreqd2_1 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_26899 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  p0enabled2 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_26903 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  p1enabled2 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {32{`RANDOM}};
  p0Datad3 = _RAND_262[1023:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  p0Validd3 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {32{`RANDOM}};
  p1Datad3 = _RAND_264[1023:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  p1Validd3 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {32{`RANDOM}};
  p2Datad3 = _RAND_266[1023:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  p2Validd3 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {32{`RANDOM}};
  _T_27292 = _RAND_268[1023:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {32{`RANDOM}};
  _T_27294 = _RAND_269[1023:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {32{`RANDOM}};
  p0Datad6 = _RAND_270[1023:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_27298 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_27300 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  p0Validd6 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {32{`RANDOM}};
  _T_27304 = _RAND_274[1023:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {32{`RANDOM}};
  _T_27306 = _RAND_275[1023:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {32{`RANDOM}};
  p1Datad6 = _RAND_276[1023:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_27310 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_27312 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  p1Validd6 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {32{`RANDOM}};
  _T_27316 = _RAND_280[1023:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {32{`RANDOM}};
  _T_27318 = _RAND_281[1023:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {32{`RANDOM}};
  p2Datad6 = _RAND_282[1023:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_27322 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_27324 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  p2Validd6 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ramWreqd1_0_0 <= 1'h0;
    end else begin
      if (4'h0 == _T_1533) begin
        ramWreqd1_0_0 <= _T_1559;
      end else begin
        ramWreqd1_0_0 <= 1'h0;
      end
    end
    if (reset) begin
      ramWreqd1_0_1 <= 1'h0;
    end else begin
      if (4'h0 == _T_1533) begin
        ramWreqd1_0_1 <= _T_1586;
      end else begin
        ramWreqd1_0_1 <= 1'h0;
      end
    end
    if (reset) begin
      ramWreqd1_1_0 <= 1'h0;
    end else begin
      ramWreqd1_1_0 <= _T_4142;
    end
    if (reset) begin
      ramWreqd1_1_1 <= 1'h0;
    end else begin
      ramWreqd1_1_1 <= _T_4143;
    end
    if (reset) begin
      ramWreqd1_2_0 <= 1'h0;
    end else begin
      ramWreqd1_2_0 <= _T_4144;
    end
    if (reset) begin
      ramWreqd1_2_1 <= 1'h0;
    end else begin
      ramWreqd1_2_1 <= _T_4145;
    end
    if (reset) begin
      ramWreqd1_3_0 <= 1'h0;
    end else begin
      ramWreqd1_3_0 <= _T_4146;
    end
    if (reset) begin
      ramWreqd1_3_1 <= 1'h0;
    end else begin
      ramWreqd1_3_1 <= _T_4147;
    end
    if (reset) begin
      ramWreqd1_4_0 <= 1'h0;
    end else begin
      ramWreqd1_4_0 <= _T_4148;
    end
    if (reset) begin
      ramWreqd1_4_1 <= 1'h0;
    end else begin
      ramWreqd1_4_1 <= _T_4149;
    end
    if (reset) begin
      ramWreqd1_5_0 <= 1'h0;
    end else begin
      ramWreqd1_5_0 <= _T_4150;
    end
    if (reset) begin
      ramWreqd1_5_1 <= 1'h0;
    end else begin
      ramWreqd1_5_1 <= _T_4151;
    end
    if (reset) begin
      ramWreqd1_6_0 <= 1'h0;
    end else begin
      ramWreqd1_6_0 <= _T_4152;
    end
    if (reset) begin
      ramWreqd1_6_1 <= 1'h0;
    end else begin
      ramWreqd1_6_1 <= _T_4153;
    end
    if (reset) begin
      ramWreqd1_7_0 <= 1'h0;
    end else begin
      ramWreqd1_7_0 <= _T_4154;
    end
    if (reset) begin
      ramWreqd1_7_1 <= 1'h0;
    end else begin
      ramWreqd1_7_1 <= _T_4155;
    end
    if (reset) begin
      ramWreqd1_8_0 <= 1'h0;
    end else begin
      ramWreqd1_8_0 <= _T_4156;
    end
    if (reset) begin
      ramWreqd1_8_1 <= 1'h0;
    end else begin
      ramWreqd1_8_1 <= _T_4157;
    end
    if (reset) begin
      ramWreqd1_9_0 <= 1'h0;
    end else begin
      ramWreqd1_9_0 <= _T_4158;
    end
    if (reset) begin
      ramWreqd1_9_1 <= 1'h0;
    end else begin
      ramWreqd1_9_1 <= _T_4159;
    end
    if (reset) begin
      ramWreqd1_10_0 <= 1'h0;
    end else begin
      ramWreqd1_10_0 <= _T_4160;
    end
    if (reset) begin
      ramWreqd1_10_1 <= 1'h0;
    end else begin
      ramWreqd1_10_1 <= _T_4161;
    end
    if (reset) begin
      ramWreqd1_11_0 <= 1'h0;
    end else begin
      ramWreqd1_11_0 <= _T_4162;
    end
    if (reset) begin
      ramWreqd1_11_1 <= 1'h0;
    end else begin
      ramWreqd1_11_1 <= _T_4163;
    end
    if (reset) begin
      ramWreqd1_12_0 <= 1'h0;
    end else begin
      ramWreqd1_12_0 <= _T_4164;
    end
    if (reset) begin
      ramWreqd1_12_1 <= 1'h0;
    end else begin
      ramWreqd1_12_1 <= _T_4165;
    end
    if (reset) begin
      ramWreqd1_13_0 <= 1'h0;
    end else begin
      ramWreqd1_13_0 <= _T_4166;
    end
    if (reset) begin
      ramWreqd1_13_1 <= 1'h0;
    end else begin
      ramWreqd1_13_1 <= _T_4167;
    end
    if (reset) begin
      ramWreqd1_14_0 <= 1'h0;
    end else begin
      ramWreqd1_14_0 <= _T_4168;
    end
    if (reset) begin
      ramWreqd1_14_1 <= 1'h0;
    end else begin
      ramWreqd1_14_1 <= _T_4169;
    end
    if (reset) begin
      ramWreqd1_15_0 <= 1'h0;
    end else begin
      if (4'hf == _T_1587) begin
        ramWreqd1_15_0 <= _T_1615;
      end else begin
        ramWreqd1_15_0 <= 1'h0;
      end
    end
    if (reset) begin
      ramWreqd1_15_1 <= 1'h0;
    end else begin
      if (4'hf == _T_1587) begin
        ramWreqd1_15_1 <= _T_1642;
      end else begin
        ramWreqd1_15_1 <= 1'h0;
      end
    end
    ramp0Addrd1 <= io_cdma2bufDat_addr[7:0];
    ramp1Addrd1 <= io_cdma2bufWt_addr[7:0];
    ramp0DatLod1 <= io_cdma2bufDat_data[511:0];
    ramp0DatHid1 <= io_cdma2bufDat_data[1023:512];
    ramp1WtLod1 <= io_cdma2bufWt_data[511:0];
    ramp1WtHid1 <= io_cdma2bufWt_data[511:0];
    if (reset) begin
      ramWreqd2_0_0 <= 1'h0;
    end else begin
      ramWreqd2_0_0 <= ramWreqd1_0_0;
    end
    if (reset) begin
      ramWreqd2_0_1 <= 1'h0;
    end else begin
      ramWreqd2_0_1 <= ramWreqd1_0_1;
    end
    if (reset) begin
      ramWreqd2_1_0 <= 1'h0;
    end else begin
      ramWreqd2_1_0 <= ramWreqd1_1_0;
    end
    if (reset) begin
      ramWreqd2_1_1 <= 1'h0;
    end else begin
      ramWreqd2_1_1 <= ramWreqd1_1_1;
    end
    if (reset) begin
      ramWreqd2_2_0 <= 1'h0;
    end else begin
      ramWreqd2_2_0 <= ramWreqd1_2_0;
    end
    if (reset) begin
      ramWreqd2_2_1 <= 1'h0;
    end else begin
      ramWreqd2_2_1 <= ramWreqd1_2_1;
    end
    if (reset) begin
      ramWreqd2_3_0 <= 1'h0;
    end else begin
      ramWreqd2_3_0 <= ramWreqd1_3_0;
    end
    if (reset) begin
      ramWreqd2_3_1 <= 1'h0;
    end else begin
      ramWreqd2_3_1 <= ramWreqd1_3_1;
    end
    if (reset) begin
      ramWreqd2_4_0 <= 1'h0;
    end else begin
      ramWreqd2_4_0 <= ramWreqd1_4_0;
    end
    if (reset) begin
      ramWreqd2_4_1 <= 1'h0;
    end else begin
      ramWreqd2_4_1 <= ramWreqd1_4_1;
    end
    if (reset) begin
      ramWreqd2_5_0 <= 1'h0;
    end else begin
      ramWreqd2_5_0 <= ramWreqd1_5_0;
    end
    if (reset) begin
      ramWreqd2_5_1 <= 1'h0;
    end else begin
      ramWreqd2_5_1 <= ramWreqd1_5_1;
    end
    if (reset) begin
      ramWreqd2_6_0 <= 1'h0;
    end else begin
      ramWreqd2_6_0 <= ramWreqd1_6_0;
    end
    if (reset) begin
      ramWreqd2_6_1 <= 1'h0;
    end else begin
      ramWreqd2_6_1 <= ramWreqd1_6_1;
    end
    if (reset) begin
      ramWreqd2_7_0 <= 1'h0;
    end else begin
      ramWreqd2_7_0 <= ramWreqd1_7_0;
    end
    if (reset) begin
      ramWreqd2_7_1 <= 1'h0;
    end else begin
      ramWreqd2_7_1 <= ramWreqd1_7_1;
    end
    if (reset) begin
      ramWreqd2_8_0 <= 1'h0;
    end else begin
      ramWreqd2_8_0 <= ramWreqd1_8_0;
    end
    if (reset) begin
      ramWreqd2_8_1 <= 1'h0;
    end else begin
      ramWreqd2_8_1 <= ramWreqd1_8_1;
    end
    if (reset) begin
      ramWreqd2_9_0 <= 1'h0;
    end else begin
      ramWreqd2_9_0 <= ramWreqd1_9_0;
    end
    if (reset) begin
      ramWreqd2_9_1 <= 1'h0;
    end else begin
      ramWreqd2_9_1 <= ramWreqd1_9_1;
    end
    if (reset) begin
      ramWreqd2_10_0 <= 1'h0;
    end else begin
      ramWreqd2_10_0 <= ramWreqd1_10_0;
    end
    if (reset) begin
      ramWreqd2_10_1 <= 1'h0;
    end else begin
      ramWreqd2_10_1 <= ramWreqd1_10_1;
    end
    if (reset) begin
      ramWreqd2_11_0 <= 1'h0;
    end else begin
      ramWreqd2_11_0 <= ramWreqd1_11_0;
    end
    if (reset) begin
      ramWreqd2_11_1 <= 1'h0;
    end else begin
      ramWreqd2_11_1 <= ramWreqd1_11_1;
    end
    if (reset) begin
      ramWreqd2_12_0 <= 1'h0;
    end else begin
      ramWreqd2_12_0 <= ramWreqd1_12_0;
    end
    if (reset) begin
      ramWreqd2_12_1 <= 1'h0;
    end else begin
      ramWreqd2_12_1 <= ramWreqd1_12_1;
    end
    if (reset) begin
      ramWreqd2_13_0 <= 1'h0;
    end else begin
      ramWreqd2_13_0 <= ramWreqd1_13_0;
    end
    if (reset) begin
      ramWreqd2_13_1 <= 1'h0;
    end else begin
      ramWreqd2_13_1 <= ramWreqd1_13_1;
    end
    if (reset) begin
      ramWreqd2_14_0 <= 1'h0;
    end else begin
      ramWreqd2_14_0 <= ramWreqd1_14_0;
    end
    if (reset) begin
      ramWreqd2_14_1 <= 1'h0;
    end else begin
      ramWreqd2_14_1 <= ramWreqd1_14_1;
    end
    if (reset) begin
      ramWreqd2_15_0 <= 1'h0;
    end else begin
      ramWreqd2_15_0 <= ramWreqd1_15_0;
    end
    if (reset) begin
      ramWreqd2_15_1 <= 1'h0;
    end else begin
      ramWreqd2_15_1 <= ramWreqd1_15_1;
    end
    if (reset) begin
      ramRreq_0_0 <= 1'h0;
    end else begin
      if (4'h0 == _T_10644) begin
        ramRreq_0_0 <= io_sc2bufDat_enable;
      end else begin
        ramRreq_0_0 <= 1'h0;
      end
    end
    if (reset) begin
      ramRreq_0_1 <= 1'h0;
    end else begin
      if (4'h0 == _T_10644) begin
        ramRreq_0_1 <= io_sc2bufDat_enable;
      end else begin
        ramRreq_0_1 <= 1'h0;
      end
    end
    if (reset) begin
      ramRreq_1_0 <= 1'h0;
    end else begin
      ramRreq_1_0 <= _T_15704;
    end
    if (reset) begin
      ramRreq_1_1 <= 1'h0;
    end else begin
      ramRreq_1_1 <= _T_15704;
    end
    if (reset) begin
      ramRreq_2_0 <= 1'h0;
    end else begin
      ramRreq_2_0 <= _T_15706;
    end
    if (reset) begin
      ramRreq_2_1 <= 1'h0;
    end else begin
      ramRreq_2_1 <= _T_15706;
    end
    if (reset) begin
      ramRreq_3_0 <= 1'h0;
    end else begin
      ramRreq_3_0 <= _T_15708;
    end
    if (reset) begin
      ramRreq_3_1 <= 1'h0;
    end else begin
      ramRreq_3_1 <= _T_15708;
    end
    if (reset) begin
      ramRreq_4_0 <= 1'h0;
    end else begin
      ramRreq_4_0 <= _T_15710;
    end
    if (reset) begin
      ramRreq_4_1 <= 1'h0;
    end else begin
      ramRreq_4_1 <= _T_15710;
    end
    if (reset) begin
      ramRreq_5_0 <= 1'h0;
    end else begin
      ramRreq_5_0 <= _T_15712;
    end
    if (reset) begin
      ramRreq_5_1 <= 1'h0;
    end else begin
      ramRreq_5_1 <= _T_15712;
    end
    if (reset) begin
      ramRreq_6_0 <= 1'h0;
    end else begin
      ramRreq_6_0 <= _T_15714;
    end
    if (reset) begin
      ramRreq_6_1 <= 1'h0;
    end else begin
      ramRreq_6_1 <= _T_15714;
    end
    if (reset) begin
      ramRreq_7_0 <= 1'h0;
    end else begin
      ramRreq_7_0 <= _T_15716;
    end
    if (reset) begin
      ramRreq_7_1 <= 1'h0;
    end else begin
      ramRreq_7_1 <= _T_15716;
    end
    if (reset) begin
      ramRreq_8_0 <= 1'h0;
    end else begin
      ramRreq_8_0 <= _T_15718;
    end
    if (reset) begin
      ramRreq_8_1 <= 1'h0;
    end else begin
      ramRreq_8_1 <= _T_15718;
    end
    if (reset) begin
      ramRreq_9_0 <= 1'h0;
    end else begin
      ramRreq_9_0 <= _T_15720;
    end
    if (reset) begin
      ramRreq_9_1 <= 1'h0;
    end else begin
      ramRreq_9_1 <= _T_15720;
    end
    if (reset) begin
      ramRreq_10_0 <= 1'h0;
    end else begin
      ramRreq_10_0 <= _T_15722;
    end
    if (reset) begin
      ramRreq_10_1 <= 1'h0;
    end else begin
      ramRreq_10_1 <= _T_15722;
    end
    if (reset) begin
      ramRreq_11_0 <= 1'h0;
    end else begin
      ramRreq_11_0 <= _T_15724;
    end
    if (reset) begin
      ramRreq_11_1 <= 1'h0;
    end else begin
      ramRreq_11_1 <= _T_15724;
    end
    if (reset) begin
      ramRreq_12_0 <= 1'h0;
    end else begin
      ramRreq_12_0 <= _T_15726;
    end
    if (reset) begin
      ramRreq_12_1 <= 1'h0;
    end else begin
      ramRreq_12_1 <= _T_15726;
    end
    if (reset) begin
      ramRreq_13_0 <= 1'h0;
    end else begin
      ramRreq_13_0 <= _T_15728;
    end
    if (reset) begin
      ramRreq_13_1 <= 1'h0;
    end else begin
      ramRreq_13_1 <= _T_15728;
    end
    if (reset) begin
      ramRreq_14_0 <= 1'h0;
    end else begin
      ramRreq_14_0 <= _T_15730;
    end
    if (reset) begin
      ramRreq_14_1 <= 1'h0;
    end else begin
      ramRreq_14_1 <= _T_15730;
    end
    if (reset) begin
      ramRreq_15_0 <= 1'h0;
    end else begin
      ramRreq_15_0 <= _T_15732;
    end
    if (reset) begin
      ramRreq_15_1 <= 1'h0;
    end else begin
      ramRreq_15_1 <= _T_15732;
    end
    if (reset) begin
      ramRaddr_0_0 <= 8'h0;
    end else begin
      ramRaddr_0_0 <= _T_15737[7:0];
    end
    if (reset) begin
      ramRaddr_0_1 <= 8'h0;
    end else begin
      ramRaddr_0_1 <= _T_15737[7:0];
    end
    if (reset) begin
      ramRaddr_1_0 <= 8'h0;
    end else begin
      ramRaddr_1_0 <= _T_15750[7:0];
    end
    if (reset) begin
      ramRaddr_1_1 <= 8'h0;
    end else begin
      ramRaddr_1_1 <= _T_15750[7:0];
    end
    if (reset) begin
      ramRaddr_2_0 <= 8'h0;
    end else begin
      ramRaddr_2_0 <= _T_15768[7:0];
    end
    if (reset) begin
      ramRaddr_2_1 <= 8'h0;
    end else begin
      ramRaddr_2_1 <= _T_15768[7:0];
    end
    if (reset) begin
      ramRaddr_3_0 <= 8'h0;
    end else begin
      ramRaddr_3_0 <= _T_15786[7:0];
    end
    if (reset) begin
      ramRaddr_3_1 <= 8'h0;
    end else begin
      ramRaddr_3_1 <= _T_15786[7:0];
    end
    if (reset) begin
      ramRaddr_4_0 <= 8'h0;
    end else begin
      ramRaddr_4_0 <= _T_15804[7:0];
    end
    if (reset) begin
      ramRaddr_4_1 <= 8'h0;
    end else begin
      ramRaddr_4_1 <= _T_15804[7:0];
    end
    if (reset) begin
      ramRaddr_5_0 <= 8'h0;
    end else begin
      ramRaddr_5_0 <= _T_15822[7:0];
    end
    if (reset) begin
      ramRaddr_5_1 <= 8'h0;
    end else begin
      ramRaddr_5_1 <= _T_15822[7:0];
    end
    if (reset) begin
      ramRaddr_6_0 <= 8'h0;
    end else begin
      ramRaddr_6_0 <= _T_15840[7:0];
    end
    if (reset) begin
      ramRaddr_6_1 <= 8'h0;
    end else begin
      ramRaddr_6_1 <= _T_15840[7:0];
    end
    if (reset) begin
      ramRaddr_7_0 <= 8'h0;
    end else begin
      ramRaddr_7_0 <= _T_15858[7:0];
    end
    if (reset) begin
      ramRaddr_7_1 <= 8'h0;
    end else begin
      ramRaddr_7_1 <= _T_15858[7:0];
    end
    if (reset) begin
      ramRaddr_8_0 <= 8'h0;
    end else begin
      ramRaddr_8_0 <= _T_15876[7:0];
    end
    if (reset) begin
      ramRaddr_8_1 <= 8'h0;
    end else begin
      ramRaddr_8_1 <= _T_15876[7:0];
    end
    if (reset) begin
      ramRaddr_9_0 <= 8'h0;
    end else begin
      ramRaddr_9_0 <= _T_15894[7:0];
    end
    if (reset) begin
      ramRaddr_9_1 <= 8'h0;
    end else begin
      ramRaddr_9_1 <= _T_15894[7:0];
    end
    if (reset) begin
      ramRaddr_10_0 <= 8'h0;
    end else begin
      ramRaddr_10_0 <= _T_15912[7:0];
    end
    if (reset) begin
      ramRaddr_10_1 <= 8'h0;
    end else begin
      ramRaddr_10_1 <= _T_15912[7:0];
    end
    if (reset) begin
      ramRaddr_11_0 <= 8'h0;
    end else begin
      ramRaddr_11_0 <= _T_15930[7:0];
    end
    if (reset) begin
      ramRaddr_11_1 <= 8'h0;
    end else begin
      ramRaddr_11_1 <= _T_15930[7:0];
    end
    if (reset) begin
      ramRaddr_12_0 <= 8'h0;
    end else begin
      ramRaddr_12_0 <= _T_15948[7:0];
    end
    if (reset) begin
      ramRaddr_12_1 <= 8'h0;
    end else begin
      ramRaddr_12_1 <= _T_15948[7:0];
    end
    if (reset) begin
      ramRaddr_13_0 <= 8'h0;
    end else begin
      ramRaddr_13_0 <= _T_15966[7:0];
    end
    if (reset) begin
      ramRaddr_13_1 <= 8'h0;
    end else begin
      ramRaddr_13_1 <= _T_15966[7:0];
    end
    if (reset) begin
      ramRaddr_14_0 <= 8'h0;
    end else begin
      ramRaddr_14_0 <= _T_15984[7:0];
    end
    if (reset) begin
      ramRaddr_14_1 <= 8'h0;
    end else begin
      ramRaddr_14_1 <= _T_15984[7:0];
    end
    if (reset) begin
      ramRaddr_15_0 <= 8'h0;
    end else begin
      ramRaddr_15_0 <= _T_16002[7:0];
    end
    if (reset) begin
      ramRaddr_15_1 <= 8'h0;
    end else begin
      ramRaddr_15_1 <= _T_16002[7:0];
    end
    if (4'h0 == _T_10644) begin
      _T_16712_0_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_0_0 <= 1'h0;
    end
    if (4'h0 == _T_10644) begin
      _T_16712_0_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_0_1 <= 1'h0;
    end
    if (4'h1 == _T_10644) begin
      _T_16712_1_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_1_0 <= 1'h0;
    end
    if (4'h1 == _T_10644) begin
      _T_16712_1_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_1_1 <= 1'h0;
    end
    if (4'h2 == _T_10644) begin
      _T_16712_2_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_2_0 <= 1'h0;
    end
    if (4'h2 == _T_10644) begin
      _T_16712_2_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_2_1 <= 1'h0;
    end
    if (4'h3 == _T_10644) begin
      _T_16712_3_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_3_0 <= 1'h0;
    end
    if (4'h3 == _T_10644) begin
      _T_16712_3_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_3_1 <= 1'h0;
    end
    if (4'h4 == _T_10644) begin
      _T_16712_4_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_4_0 <= 1'h0;
    end
    if (4'h4 == _T_10644) begin
      _T_16712_4_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_4_1 <= 1'h0;
    end
    if (4'h5 == _T_10644) begin
      _T_16712_5_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_5_0 <= 1'h0;
    end
    if (4'h5 == _T_10644) begin
      _T_16712_5_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_5_1 <= 1'h0;
    end
    if (4'h6 == _T_10644) begin
      _T_16712_6_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_6_0 <= 1'h0;
    end
    if (4'h6 == _T_10644) begin
      _T_16712_6_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_6_1 <= 1'h0;
    end
    if (4'h7 == _T_10644) begin
      _T_16712_7_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_7_0 <= 1'h0;
    end
    if (4'h7 == _T_10644) begin
      _T_16712_7_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_7_1 <= 1'h0;
    end
    if (4'h8 == _T_10644) begin
      _T_16712_8_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_8_0 <= 1'h0;
    end
    if (4'h8 == _T_10644) begin
      _T_16712_8_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_8_1 <= 1'h0;
    end
    if (4'h9 == _T_10644) begin
      _T_16712_9_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_9_0 <= 1'h0;
    end
    if (4'h9 == _T_10644) begin
      _T_16712_9_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_9_1 <= 1'h0;
    end
    if (4'ha == _T_10644) begin
      _T_16712_10_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_10_0 <= 1'h0;
    end
    if (4'ha == _T_10644) begin
      _T_16712_10_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_10_1 <= 1'h0;
    end
    if (4'hb == _T_10644) begin
      _T_16712_11_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_11_0 <= 1'h0;
    end
    if (4'hb == _T_10644) begin
      _T_16712_11_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_11_1 <= 1'h0;
    end
    if (4'hc == _T_10644) begin
      _T_16712_12_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_12_0 <= 1'h0;
    end
    if (4'hc == _T_10644) begin
      _T_16712_12_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_12_1 <= 1'h0;
    end
    if (4'hd == _T_10644) begin
      _T_16712_13_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_13_0 <= 1'h0;
    end
    if (4'hd == _T_10644) begin
      _T_16712_13_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_13_1 <= 1'h0;
    end
    if (4'he == _T_10644) begin
      _T_16712_14_0 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_14_0 <= 1'h0;
    end
    if (4'he == _T_10644) begin
      _T_16712_14_1 <= io_sc2bufDat_enable;
    end else begin
      _T_16712_14_1 <= 1'h0;
    end
    datRreqd2_0_0 <= _T_16712_0_0;
    datRreqd2_0_1 <= _T_16712_0_1;
    datRreqd2_1_0 <= _T_16712_1_0;
    datRreqd2_1_1 <= _T_16712_1_1;
    datRreqd2_2_0 <= _T_16712_2_0;
    datRreqd2_2_1 <= _T_16712_2_1;
    datRreqd2_3_0 <= _T_16712_3_0;
    datRreqd2_3_1 <= _T_16712_3_1;
    datRreqd2_4_0 <= _T_16712_4_0;
    datRreqd2_4_1 <= _T_16712_4_1;
    datRreqd2_5_0 <= _T_16712_5_0;
    datRreqd2_5_1 <= _T_16712_5_1;
    datRreqd2_6_0 <= _T_16712_6_0;
    datRreqd2_6_1 <= _T_16712_6_1;
    datRreqd2_7_0 <= _T_16712_7_0;
    datRreqd2_7_1 <= _T_16712_7_1;
    datRreqd2_8_0 <= _T_16712_8_0;
    datRreqd2_8_1 <= _T_16712_8_1;
    datRreqd2_9_0 <= _T_16712_9_0;
    datRreqd2_9_1 <= _T_16712_9_1;
    datRreqd2_10_0 <= _T_16712_10_0;
    datRreqd2_10_1 <= _T_16712_10_1;
    datRreqd2_11_0 <= _T_16712_11_0;
    datRreqd2_11_1 <= _T_16712_11_1;
    datRreqd2_12_0 <= _T_16712_12_0;
    datRreqd2_12_1 <= _T_16712_12_1;
    datRreqd2_13_0 <= _T_16712_13_0;
    datRreqd2_13_1 <= _T_16712_13_1;
    datRreqd2_14_0 <= _T_16712_14_0;
    datRreqd2_14_1 <= _T_16712_14_1;
    if (4'h1 == _T_10687) begin
      _T_21752_1_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_1_0 <= 1'h0;
    end
    if (4'h1 == _T_10687) begin
      _T_21752_1_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_1_1 <= 1'h0;
    end
    if (4'h2 == _T_10687) begin
      _T_21752_2_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_2_0 <= 1'h0;
    end
    if (4'h2 == _T_10687) begin
      _T_21752_2_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_2_1 <= 1'h0;
    end
    if (4'h3 == _T_10687) begin
      _T_21752_3_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_3_0 <= 1'h0;
    end
    if (4'h3 == _T_10687) begin
      _T_21752_3_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_3_1 <= 1'h0;
    end
    if (4'h4 == _T_10687) begin
      _T_21752_4_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_4_0 <= 1'h0;
    end
    if (4'h4 == _T_10687) begin
      _T_21752_4_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_4_1 <= 1'h0;
    end
    if (4'h5 == _T_10687) begin
      _T_21752_5_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_5_0 <= 1'h0;
    end
    if (4'h5 == _T_10687) begin
      _T_21752_5_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_5_1 <= 1'h0;
    end
    if (4'h6 == _T_10687) begin
      _T_21752_6_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_6_0 <= 1'h0;
    end
    if (4'h6 == _T_10687) begin
      _T_21752_6_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_6_1 <= 1'h0;
    end
    if (4'h7 == _T_10687) begin
      _T_21752_7_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_7_0 <= 1'h0;
    end
    if (4'h7 == _T_10687) begin
      _T_21752_7_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_7_1 <= 1'h0;
    end
    if (4'h8 == _T_10687) begin
      _T_21752_8_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_8_0 <= 1'h0;
    end
    if (4'h8 == _T_10687) begin
      _T_21752_8_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_8_1 <= 1'h0;
    end
    if (4'h9 == _T_10687) begin
      _T_21752_9_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_9_0 <= 1'h0;
    end
    if (4'h9 == _T_10687) begin
      _T_21752_9_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_9_1 <= 1'h0;
    end
    if (4'ha == _T_10687) begin
      _T_21752_10_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_10_0 <= 1'h0;
    end
    if (4'ha == _T_10687) begin
      _T_21752_10_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_10_1 <= 1'h0;
    end
    if (4'hb == _T_10687) begin
      _T_21752_11_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_11_0 <= 1'h0;
    end
    if (4'hb == _T_10687) begin
      _T_21752_11_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_11_1 <= 1'h0;
    end
    if (4'hc == _T_10687) begin
      _T_21752_12_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_12_0 <= 1'h0;
    end
    if (4'hc == _T_10687) begin
      _T_21752_12_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_12_1 <= 1'h0;
    end
    if (4'hd == _T_10687) begin
      _T_21752_13_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_13_0 <= 1'h0;
    end
    if (4'hd == _T_10687) begin
      _T_21752_13_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_13_1 <= 1'h0;
    end
    if (4'he == _T_10687) begin
      _T_21752_14_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_14_0 <= 1'h0;
    end
    if (4'he == _T_10687) begin
      _T_21752_14_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_14_1 <= 1'h0;
    end
    if (4'hf == _T_10687) begin
      _T_21752_15_0 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_15_0 <= 1'h0;
    end
    if (4'hf == _T_10687) begin
      _T_21752_15_1 <= io_sc2bufWt_enable;
    end else begin
      _T_21752_15_1 <= 1'h0;
    end
    wtRreqd2_1_0 <= _T_21752_1_0;
    wtRreqd2_1_1 <= _T_21752_1_1;
    wtRreqd2_2_0 <= _T_21752_2_0;
    wtRreqd2_2_1 <= _T_21752_2_1;
    wtRreqd2_3_0 <= _T_21752_3_0;
    wtRreqd2_3_1 <= _T_21752_3_1;
    wtRreqd2_4_0 <= _T_21752_4_0;
    wtRreqd2_4_1 <= _T_21752_4_1;
    wtRreqd2_5_0 <= _T_21752_5_0;
    wtRreqd2_5_1 <= _T_21752_5_1;
    wtRreqd2_6_0 <= _T_21752_6_0;
    wtRreqd2_6_1 <= _T_21752_6_1;
    wtRreqd2_7_0 <= _T_21752_7_0;
    wtRreqd2_7_1 <= _T_21752_7_1;
    wtRreqd2_8_0 <= _T_21752_8_0;
    wtRreqd2_8_1 <= _T_21752_8_1;
    wtRreqd2_9_0 <= _T_21752_9_0;
    wtRreqd2_9_1 <= _T_21752_9_1;
    wtRreqd2_10_0 <= _T_21752_10_0;
    wtRreqd2_10_1 <= _T_21752_10_1;
    wtRreqd2_11_0 <= _T_21752_11_0;
    wtRreqd2_11_1 <= _T_21752_11_1;
    wtRreqd2_12_0 <= _T_21752_12_0;
    wtRreqd2_12_1 <= _T_21752_12_1;
    wtRreqd2_13_0 <= _T_21752_13_0;
    wtRreqd2_13_1 <= _T_21752_13_1;
    wtRreqd2_14_0 <= _T_21752_14_0;
    wtRreqd2_14_1 <= _T_21752_14_1;
    wtRreqd2_15_0 <= _T_21752_15_0;
    wtRreqd2_15_1 <= _T_21752_15_1;
    _T_26101_0 <= io_sc2bufWMB_enable;
    _T_26101_1 <= io_sc2bufWMB_enable;
    wmbRreqd2_0 <= _T_26101_0;
    wmbRreqd2_1 <= _T_26101_1;
    _T_26899 <= io_sc2bufDat_enable;
    p0enabled2 <= _T_26899;
    _T_26903 <= io_sc2bufWt_enable;
    p1enabled2 <= _T_26903;
    p0Datad3 <= _T_27086 | _T_27073;
    p0Validd3 <= p0enabled2;
    p1Datad3 <= _T_27269 | _T_27256;
    p1Validd3 <= p1enabled2;
    p2Datad3 <= _T_27283 & _T_27255;
    p2Validd3 <= p1enabled2;
    _T_27292 <= p0Datad3;
    _T_27294 <= _T_27292;
    p0Datad6 <= _T_27294;
    _T_27298 <= p0Validd3;
    _T_27300 <= _T_27298;
    p0Validd6 <= _T_27300;
    _T_27304 <= p1Datad3;
    _T_27306 <= _T_27304;
    p1Datad6 <= _T_27306;
    _T_27310 <= p1Validd3;
    _T_27312 <= _T_27310;
    p1Validd6 <= _T_27312;
    _T_27316 <= p2Datad3;
    _T_27318 <= _T_27316;
    p2Datad6 <= _T_27318;
    _T_27322 <= p2Validd3;
    _T_27324 <= _T_27322;
    p2Validd6 <= _T_27324;
  end
endmodule
