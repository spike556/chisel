module FMul( // @[:@3.2]
  input  [162:0] io_a, // @[:@6.4]
  input  [15:0]  io_b, // @[:@6.4]
  output [177:0] io_pout // @[:@6.4]
);
  wire  _T_84; // @[PEAlter.scala 19:15:@60.4]
  wire [163:0] _GEN_16; // @[PEAlter.scala 20:34:@63.6]
  wire [163:0] _T_88; // @[PEAlter.scala 20:34:@63.6]
  wire [177:0] _T_89; // @[PEAlter.scala 20:26:@64.6]
  wire [177:0] tmp_1; // @[PEAlter.scala 19:28:@62.4]
  wire  _T_90; // @[PEAlter.scala 19:15:@70.4]
  wire [163:0] _T_94; // @[PEAlter.scala 20:34:@73.6]
  wire [177:0] _GEN_18; // @[PEAlter.scala 20:26:@74.6]
  wire [177:0] _T_95; // @[PEAlter.scala 20:26:@74.6]
  wire [177:0] tmp_2; // @[PEAlter.scala 19:28:@72.4]
  wire  _T_96; // @[PEAlter.scala 19:15:@80.4]
  wire [165:0] _GEN_19; // @[PEAlter.scala 20:34:@83.6]
  wire [165:0] _T_100; // @[PEAlter.scala 20:34:@83.6]
  wire [177:0] _GEN_20; // @[PEAlter.scala 20:26:@84.6]
  wire [177:0] _T_101; // @[PEAlter.scala 20:26:@84.6]
  wire [177:0] tmp_3; // @[PEAlter.scala 19:28:@82.4]
  wire  _T_102; // @[PEAlter.scala 19:15:@90.4]
  wire [165:0] _T_106; // @[PEAlter.scala 20:34:@93.6]
  wire [177:0] _GEN_22; // @[PEAlter.scala 20:26:@94.6]
  wire [177:0] _T_107; // @[PEAlter.scala 20:26:@94.6]
  wire [177:0] tmp_4; // @[PEAlter.scala 19:28:@92.4]
  wire  _T_108; // @[PEAlter.scala 19:15:@100.4]
  wire [169:0] _GEN_23; // @[PEAlter.scala 20:34:@103.6]
  wire [169:0] _T_112; // @[PEAlter.scala 20:34:@103.6]
  wire [177:0] _GEN_24; // @[PEAlter.scala 20:26:@104.6]
  wire [177:0] _T_113; // @[PEAlter.scala 20:26:@104.6]
  wire [177:0] tmp_5; // @[PEAlter.scala 19:28:@102.4]
  wire  _T_114; // @[PEAlter.scala 19:15:@110.4]
  wire [169:0] _T_118; // @[PEAlter.scala 20:34:@113.6]
  wire [177:0] _GEN_26; // @[PEAlter.scala 20:26:@114.6]
  wire [177:0] _T_119; // @[PEAlter.scala 20:26:@114.6]
  wire [177:0] tmp_6; // @[PEAlter.scala 19:28:@112.4]
  wire  _T_120; // @[PEAlter.scala 19:15:@120.4]
  wire [169:0] _T_124; // @[PEAlter.scala 20:34:@123.6]
  wire [177:0] _GEN_28; // @[PEAlter.scala 20:26:@124.6]
  wire [177:0] _T_125; // @[PEAlter.scala 20:26:@124.6]
  wire [177:0] tmp_7; // @[PEAlter.scala 19:28:@122.4]
  wire  _T_126; // @[PEAlter.scala 19:15:@130.4]
  wire [169:0] _T_130; // @[PEAlter.scala 20:34:@133.6]
  wire [177:0] _GEN_30; // @[PEAlter.scala 20:26:@134.6]
  wire [177:0] _T_131; // @[PEAlter.scala 20:26:@134.6]
  wire [177:0] tmp_8; // @[PEAlter.scala 19:28:@132.4]
  wire  _T_132; // @[PEAlter.scala 19:15:@140.4]
  wire [177:0] _GEN_31; // @[PEAlter.scala 20:34:@143.6]
  wire [177:0] _T_136; // @[PEAlter.scala 20:34:@143.6]
  wire [177:0] _T_137; // @[PEAlter.scala 20:26:@144.6]
  wire [177:0] tmp_9; // @[PEAlter.scala 19:28:@142.4]
  wire  _T_138; // @[PEAlter.scala 19:15:@150.4]
  wire [177:0] _T_142; // @[PEAlter.scala 20:34:@153.6]
  wire [177:0] _T_143; // @[PEAlter.scala 20:26:@154.6]
  wire [177:0] tmp_10; // @[PEAlter.scala 19:28:@152.4]
  wire  _T_144; // @[PEAlter.scala 19:15:@160.4]
  wire [177:0] _T_148; // @[PEAlter.scala 20:34:@163.6]
  wire [177:0] _T_149; // @[PEAlter.scala 20:26:@164.6]
  wire [177:0] tmp_11; // @[PEAlter.scala 19:28:@162.4]
  wire  _T_150; // @[PEAlter.scala 19:15:@170.4]
  wire [177:0] _T_154; // @[PEAlter.scala 20:34:@173.6]
  wire [177:0] _T_155; // @[PEAlter.scala 20:26:@174.6]
  wire [177:0] tmp_12; // @[PEAlter.scala 19:28:@172.4]
  wire  _T_156; // @[PEAlter.scala 19:15:@180.4]
  wire [177:0] _T_160; // @[PEAlter.scala 20:34:@183.6]
  wire [177:0] _T_161; // @[PEAlter.scala 20:26:@184.6]
  wire [177:0] tmp_13; // @[PEAlter.scala 19:28:@182.4]
  wire  _T_162; // @[PEAlter.scala 19:15:@190.4]
  wire [177:0] _T_166; // @[PEAlter.scala 20:34:@193.6]
  wire [177:0] _T_167; // @[PEAlter.scala 20:26:@194.6]
  wire [177:0] tmp_14; // @[PEAlter.scala 19:28:@192.4]
  wire  _T_168; // @[PEAlter.scala 19:15:@200.4]
  wire [177:0] _T_172; // @[PEAlter.scala 20:34:@203.6]
  wire [177:0] _T_173; // @[PEAlter.scala 20:26:@204.6]
  wire [177:0] tmp_15; // @[PEAlter.scala 19:28:@202.4]
  wire  _T_174; // @[PEAlter.scala 19:15:@210.4]
  wire [177:0] _T_178; // @[PEAlter.scala 20:34:@213.6]
  wire [177:0] _T_179; // @[PEAlter.scala 20:26:@214.6]
  assign _T_84 = io_b[0]; // @[PEAlter.scala 19:15:@60.4]
  assign _GEN_16 = {{1'd0}, io_a}; // @[PEAlter.scala 20:34:@63.6]
  assign _T_88 = _GEN_16 << 1'h0; // @[PEAlter.scala 20:34:@63.6]
  assign _T_89 = {{14'd0}, _T_88}; // @[PEAlter.scala 20:26:@64.6]
  assign tmp_1 = _T_84 ? _T_89 : 178'h0; // @[PEAlter.scala 19:28:@62.4]
  assign _T_90 = io_b[1]; // @[PEAlter.scala 19:15:@70.4]
  assign _T_94 = _GEN_16 << 1'h1; // @[PEAlter.scala 20:34:@73.6]
  assign _GEN_18 = {{14'd0}, _T_94}; // @[PEAlter.scala 20:26:@74.6]
  assign _T_95 = tmp_1 ^ _GEN_18; // @[PEAlter.scala 20:26:@74.6]
  assign tmp_2 = _T_90 ? _T_95 : tmp_1; // @[PEAlter.scala 19:28:@72.4]
  assign _T_96 = io_b[2]; // @[PEAlter.scala 19:15:@80.4]
  assign _GEN_19 = {{3'd0}, io_a}; // @[PEAlter.scala 20:34:@83.6]
  assign _T_100 = _GEN_19 << 2'h2; // @[PEAlter.scala 20:34:@83.6]
  assign _GEN_20 = {{12'd0}, _T_100}; // @[PEAlter.scala 20:26:@84.6]
  assign _T_101 = tmp_2 ^ _GEN_20; // @[PEAlter.scala 20:26:@84.6]
  assign tmp_3 = _T_96 ? _T_101 : tmp_2; // @[PEAlter.scala 19:28:@82.4]
  assign _T_102 = io_b[3]; // @[PEAlter.scala 19:15:@90.4]
  assign _T_106 = _GEN_19 << 2'h3; // @[PEAlter.scala 20:34:@93.6]
  assign _GEN_22 = {{12'd0}, _T_106}; // @[PEAlter.scala 20:26:@94.6]
  assign _T_107 = tmp_3 ^ _GEN_22; // @[PEAlter.scala 20:26:@94.6]
  assign tmp_4 = _T_102 ? _T_107 : tmp_3; // @[PEAlter.scala 19:28:@92.4]
  assign _T_108 = io_b[4]; // @[PEAlter.scala 19:15:@100.4]
  assign _GEN_23 = {{7'd0}, io_a}; // @[PEAlter.scala 20:34:@103.6]
  assign _T_112 = _GEN_23 << 3'h4; // @[PEAlter.scala 20:34:@103.6]
  assign _GEN_24 = {{8'd0}, _T_112}; // @[PEAlter.scala 20:26:@104.6]
  assign _T_113 = tmp_4 ^ _GEN_24; // @[PEAlter.scala 20:26:@104.6]
  assign tmp_5 = _T_108 ? _T_113 : tmp_4; // @[PEAlter.scala 19:28:@102.4]
  assign _T_114 = io_b[5]; // @[PEAlter.scala 19:15:@110.4]
  assign _T_118 = _GEN_23 << 3'h5; // @[PEAlter.scala 20:34:@113.6]
  assign _GEN_26 = {{8'd0}, _T_118}; // @[PEAlter.scala 20:26:@114.6]
  assign _T_119 = tmp_5 ^ _GEN_26; // @[PEAlter.scala 20:26:@114.6]
  assign tmp_6 = _T_114 ? _T_119 : tmp_5; // @[PEAlter.scala 19:28:@112.4]
  assign _T_120 = io_b[6]; // @[PEAlter.scala 19:15:@120.4]
  assign _T_124 = _GEN_23 << 3'h6; // @[PEAlter.scala 20:34:@123.6]
  assign _GEN_28 = {{8'd0}, _T_124}; // @[PEAlter.scala 20:26:@124.6]
  assign _T_125 = tmp_6 ^ _GEN_28; // @[PEAlter.scala 20:26:@124.6]
  assign tmp_7 = _T_120 ? _T_125 : tmp_6; // @[PEAlter.scala 19:28:@122.4]
  assign _T_126 = io_b[7]; // @[PEAlter.scala 19:15:@130.4]
  assign _T_130 = _GEN_23 << 3'h7; // @[PEAlter.scala 20:34:@133.6]
  assign _GEN_30 = {{8'd0}, _T_130}; // @[PEAlter.scala 20:26:@134.6]
  assign _T_131 = tmp_7 ^ _GEN_30; // @[PEAlter.scala 20:26:@134.6]
  assign tmp_8 = _T_126 ? _T_131 : tmp_7; // @[PEAlter.scala 19:28:@132.4]
  assign _T_132 = io_b[8]; // @[PEAlter.scala 19:15:@140.4]
  assign _GEN_31 = {{15'd0}, io_a}; // @[PEAlter.scala 20:34:@143.6]
  assign _T_136 = _GEN_31 << 4'h8; // @[PEAlter.scala 20:34:@143.6]
  assign _T_137 = tmp_8 ^ _T_136; // @[PEAlter.scala 20:26:@144.6]
  assign tmp_9 = _T_132 ? _T_137 : tmp_8; // @[PEAlter.scala 19:28:@142.4]
  assign _T_138 = io_b[9]; // @[PEAlter.scala 19:15:@150.4]
  assign _T_142 = _GEN_31 << 4'h9; // @[PEAlter.scala 20:34:@153.6]
  assign _T_143 = tmp_9 ^ _T_142; // @[PEAlter.scala 20:26:@154.6]
  assign tmp_10 = _T_138 ? _T_143 : tmp_9; // @[PEAlter.scala 19:28:@152.4]
  assign _T_144 = io_b[10]; // @[PEAlter.scala 19:15:@160.4]
  assign _T_148 = _GEN_31 << 4'ha; // @[PEAlter.scala 20:34:@163.6]
  assign _T_149 = tmp_10 ^ _T_148; // @[PEAlter.scala 20:26:@164.6]
  assign tmp_11 = _T_144 ? _T_149 : tmp_10; // @[PEAlter.scala 19:28:@162.4]
  assign _T_150 = io_b[11]; // @[PEAlter.scala 19:15:@170.4]
  assign _T_154 = _GEN_31 << 4'hb; // @[PEAlter.scala 20:34:@173.6]
  assign _T_155 = tmp_11 ^ _T_154; // @[PEAlter.scala 20:26:@174.6]
  assign tmp_12 = _T_150 ? _T_155 : tmp_11; // @[PEAlter.scala 19:28:@172.4]
  assign _T_156 = io_b[12]; // @[PEAlter.scala 19:15:@180.4]
  assign _T_160 = _GEN_31 << 4'hc; // @[PEAlter.scala 20:34:@183.6]
  assign _T_161 = tmp_12 ^ _T_160; // @[PEAlter.scala 20:26:@184.6]
  assign tmp_13 = _T_156 ? _T_161 : tmp_12; // @[PEAlter.scala 19:28:@182.4]
  assign _T_162 = io_b[13]; // @[PEAlter.scala 19:15:@190.4]
  assign _T_166 = _GEN_31 << 4'hd; // @[PEAlter.scala 20:34:@193.6]
  assign _T_167 = tmp_13 ^ _T_166; // @[PEAlter.scala 20:26:@194.6]
  assign tmp_14 = _T_162 ? _T_167 : tmp_13; // @[PEAlter.scala 19:28:@192.4]
  assign _T_168 = io_b[14]; // @[PEAlter.scala 19:15:@200.4]
  assign _T_172 = _GEN_31 << 4'he; // @[PEAlter.scala 20:34:@203.6]
  assign _T_173 = tmp_14 ^ _T_172; // @[PEAlter.scala 20:26:@204.6]
  assign tmp_15 = _T_168 ? _T_173 : tmp_14; // @[PEAlter.scala 19:28:@202.4]
  assign _T_174 = io_b[15]; // @[PEAlter.scala 19:15:@210.4]
  assign _T_178 = _GEN_31 << 4'hf; // @[PEAlter.scala 20:34:@213.6]
  assign _T_179 = tmp_15 ^ _T_178; // @[PEAlter.scala 20:26:@214.6]
  assign io_pout = _T_174 ? _T_179 : tmp_15; // @[PEAlter.scala 25:11:@220.4]
endmodule
module PEAlter( // @[:@222.2]
  input          clock, // @[:@223.4]
  input  [162:0] io_a, // @[:@225.4]
  input  [162:0] io_p, // @[:@225.4]
  input  [15:0]  io_bi, // @[:@225.4]
  output [162:0] io_aout, // @[:@225.4]
  output [162:0] io_pout // @[:@225.4]
);
  wire [162:0] FMul_io_a; // @[PEAlter.scala 30:19:@228.4]
  wire [15:0] FMul_io_b; // @[PEAlter.scala 30:19:@228.4]
  wire [177:0] FMul_io_pout; // @[PEAlter.scala 30:19:@228.4]
  wire [193:0] _GEN_0; // @[PEAlter.scala 45:21:@227.4]
  wire [193:0] _T_16; // @[PEAlter.scala 45:21:@227.4]
  wire [193:0] _GEN_1; // @[PEAlter.scala 45:36:@233.4]
  wire [193:0] ptmp1; // @[PEAlter.scala 45:36:@233.4]
  wire [193:0] pGuess; // @[PEAlter.scala 46:22:@234.4]
  wire [162:0] _T_18; // @[PEAlter.scala 47:20:@235.4]
  wire [200:0] _GEN_2; // @[PEAlter.scala 47:39:@236.4]
  wire [200:0] _T_20; // @[PEAlter.scala 47:39:@236.4]
  wire [200:0] _T_22; // @[PEAlter.scala 47:57:@237.4]
  wire [200:0] _T_23; // @[PEAlter.scala 47:47:@238.4]
  wire [196:0] _GEN_4; // @[PEAlter.scala 47:75:@239.4]
  wire [196:0] _T_25; // @[PEAlter.scala 47:75:@239.4]
  wire [200:0] _GEN_5; // @[PEAlter.scala 47:65:@240.4]
  wire [200:0] _T_26; // @[PEAlter.scala 47:65:@240.4]
  wire [200:0] _T_27; // @[PEAlter.scala 47:83:@241.4]
  wire [200:0] _GEN_7; // @[PEAlter.scala 47:28:@242.4]
  reg [162:0] _T_29; // @[PEAlter.scala 50:21:@243.4]
  reg [191:0] _RAND_0;
  reg [200:0] _T_31; // @[PEAlter.scala 51:21:@246.4]
  reg [223:0] _RAND_1;
  FMul FMul ( // @[PEAlter.scala 30:19:@228.4]
    .io_a(FMul_io_a),
    .io_b(FMul_io_b),
    .io_pout(FMul_io_pout)
  );
  assign _GEN_0 = {{31'd0}, io_p}; // @[PEAlter.scala 45:21:@227.4]
  assign _T_16 = _GEN_0 << 5'h10; // @[PEAlter.scala 45:21:@227.4]
  assign _GEN_1 = {{16'd0}, FMul_io_pout}; // @[PEAlter.scala 45:36:@233.4]
  assign ptmp1 = _T_16 ^ _GEN_1; // @[PEAlter.scala 45:36:@233.4]
  assign pGuess = ptmp1 >> 8'ha3; // @[PEAlter.scala 46:22:@234.4]
  assign _T_18 = ptmp1[162:0]; // @[PEAlter.scala 47:20:@235.4]
  assign _GEN_2 = {{7'd0}, pGuess}; // @[PEAlter.scala 47:39:@236.4]
  assign _T_20 = _GEN_2 << 3'h7; // @[PEAlter.scala 47:39:@236.4]
  assign _T_22 = _GEN_2 << 3'h6; // @[PEAlter.scala 47:57:@237.4]
  assign _T_23 = _T_20 ^ _T_22; // @[PEAlter.scala 47:47:@238.4]
  assign _GEN_4 = {{3'd0}, pGuess}; // @[PEAlter.scala 47:75:@239.4]
  assign _T_25 = _GEN_4 << 2'h3; // @[PEAlter.scala 47:75:@239.4]
  assign _GEN_5 = {{4'd0}, _T_25}; // @[PEAlter.scala 47:65:@240.4]
  assign _T_26 = _T_23 ^ _GEN_5; // @[PEAlter.scala 47:65:@240.4]
  assign _T_27 = _T_26 ^ _GEN_2; // @[PEAlter.scala 47:83:@241.4]
  assign _GEN_7 = {{38'd0}, _T_18}; // @[PEAlter.scala 47:28:@242.4]
  assign io_aout = _T_29; // @[PEAlter.scala 50:11:@245.4]
  assign io_pout = _T_31[162:0]; // @[PEAlter.scala 51:11:@248.4]
  assign FMul_io_a = io_a; // @[PEAlter.scala 31:12:@231.4]
  assign FMul_io_b = io_bi; // @[PEAlter.scala 32:12:@232.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {6{`RANDOM}};
  _T_29 = _RAND_0[162:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {7{`RANDOM}};
  _T_31 = _RAND_1[200:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    _T_29 <= io_a;
    _T_31 <= _GEN_7 ^ _T_27;
  end
endmodule
module ShiftRegs( // @[:@2720.2]
  input         clock, // @[:@2721.4]
  input         reset, // @[:@2722.4]
  input  [15:0] io_in, // @[:@2723.4]
  output [15:0] io_out // @[:@2723.4]
);
  reg [15:0] delays_0; // @[ShiftRegs.scala 15:23:@2727.4]
  reg [31:0] _RAND_0;
  assign io_out = delays_0; // @[ShiftRegs.scala 24:10:@2729.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delays_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      delays_0 <= 16'h0;
    end else begin
      delays_0 <= io_in;
    end
  end
endmodule
module ShiftRegs_1( // @[:@2731.2]
  input         clock, // @[:@2732.4]
  input         reset, // @[:@2733.4]
  input  [15:0] io_in, // @[:@2734.4]
  output [15:0] io_out // @[:@2734.4]
);
  reg [15:0] delays_0; // @[ShiftRegs.scala 15:23:@2739.4]
  reg [31:0] _RAND_0;
  reg [15:0] delays_1; // @[ShiftRegs.scala 15:23:@2739.4]
  reg [31:0] _RAND_1;
  assign io_out = delays_1; // @[ShiftRegs.scala 24:10:@2742.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delays_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  delays_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      delays_0 <= 16'h0;
    end else begin
      delays_0 <= io_in;
    end
    if (reset) begin
      delays_1 <= 16'h0;
    end else begin
      delays_1 <= delays_0;
    end
  end
endmodule
module ShiftRegs_2( // @[:@2744.2]
  input         clock, // @[:@2745.4]
  input         reset, // @[:@2746.4]
  input  [15:0] io_in, // @[:@2747.4]
  output [15:0] io_out // @[:@2747.4]
);
  reg [15:0] delays_0; // @[ShiftRegs.scala 15:23:@2753.4]
  reg [31:0] _RAND_0;
  reg [15:0] delays_1; // @[ShiftRegs.scala 15:23:@2753.4]
  reg [31:0] _RAND_1;
  reg [15:0] delays_2; // @[ShiftRegs.scala 15:23:@2753.4]
  reg [31:0] _RAND_2;
  assign io_out = delays_2; // @[ShiftRegs.scala 24:10:@2757.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delays_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  delays_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delays_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      delays_0 <= 16'h0;
    end else begin
      delays_0 <= io_in;
    end
    if (reset) begin
      delays_1 <= 16'h0;
    end else begin
      delays_1 <= delays_0;
    end
    if (reset) begin
      delays_2 <= 16'h0;
    end else begin
      delays_2 <= delays_1;
    end
  end
endmodule
module ShiftRegs_3( // @[:@2759.2]
  input         clock, // @[:@2760.4]
  input         reset, // @[:@2761.4]
  input  [15:0] io_in, // @[:@2762.4]
  output [15:0] io_out // @[:@2762.4]
);
  reg [15:0] delays_0; // @[ShiftRegs.scala 15:23:@2769.4]
  reg [31:0] _RAND_0;
  reg [15:0] delays_1; // @[ShiftRegs.scala 15:23:@2769.4]
  reg [31:0] _RAND_1;
  reg [15:0] delays_2; // @[ShiftRegs.scala 15:23:@2769.4]
  reg [31:0] _RAND_2;
  reg [15:0] delays_3; // @[ShiftRegs.scala 15:23:@2769.4]
  reg [31:0] _RAND_3;
  assign io_out = delays_3; // @[ShiftRegs.scala 24:10:@2774.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delays_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  delays_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delays_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  delays_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      delays_0 <= 16'h0;
    end else begin
      delays_0 <= io_in;
    end
    if (reset) begin
      delays_1 <= 16'h0;
    end else begin
      delays_1 <= delays_0;
    end
    if (reset) begin
      delays_2 <= 16'h0;
    end else begin
      delays_2 <= delays_1;
    end
    if (reset) begin
      delays_3 <= 16'h0;
    end else begin
      delays_3 <= delays_2;
    end
  end
endmodule
module ShiftRegs_4( // @[:@2776.2]
  input         clock, // @[:@2777.4]
  input         reset, // @[:@2778.4]
  input  [15:0] io_in, // @[:@2779.4]
  output [15:0] io_out // @[:@2779.4]
);
  reg [15:0] delays_0; // @[ShiftRegs.scala 15:23:@2787.4]
  reg [31:0] _RAND_0;
  reg [15:0] delays_1; // @[ShiftRegs.scala 15:23:@2787.4]
  reg [31:0] _RAND_1;
  reg [15:0] delays_2; // @[ShiftRegs.scala 15:23:@2787.4]
  reg [31:0] _RAND_2;
  reg [15:0] delays_3; // @[ShiftRegs.scala 15:23:@2787.4]
  reg [31:0] _RAND_3;
  reg [15:0] delays_4; // @[ShiftRegs.scala 15:23:@2787.4]
  reg [31:0] _RAND_4;
  assign io_out = delays_4; // @[ShiftRegs.scala 24:10:@2793.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delays_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  delays_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delays_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  delays_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  delays_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      delays_0 <= 16'h0;
    end else begin
      delays_0 <= io_in;
    end
    if (reset) begin
      delays_1 <= 16'h0;
    end else begin
      delays_1 <= delays_0;
    end
    if (reset) begin
      delays_2 <= 16'h0;
    end else begin
      delays_2 <= delays_1;
    end
    if (reset) begin
      delays_3 <= 16'h0;
    end else begin
      delays_3 <= delays_2;
    end
    if (reset) begin
      delays_4 <= 16'h0;
    end else begin
      delays_4 <= delays_3;
    end
  end
endmodule
module ShiftRegs_5( // @[:@2795.2]
  input         clock, // @[:@2796.4]
  input         reset, // @[:@2797.4]
  input  [15:0] io_in, // @[:@2798.4]
  output [15:0] io_out // @[:@2798.4]
);
  reg [15:0] delays_0; // @[ShiftRegs.scala 15:23:@2807.4]
  reg [31:0] _RAND_0;
  reg [15:0] delays_1; // @[ShiftRegs.scala 15:23:@2807.4]
  reg [31:0] _RAND_1;
  reg [15:0] delays_2; // @[ShiftRegs.scala 15:23:@2807.4]
  reg [31:0] _RAND_2;
  reg [15:0] delays_3; // @[ShiftRegs.scala 15:23:@2807.4]
  reg [31:0] _RAND_3;
  reg [15:0] delays_4; // @[ShiftRegs.scala 15:23:@2807.4]
  reg [31:0] _RAND_4;
  reg [15:0] delays_5; // @[ShiftRegs.scala 15:23:@2807.4]
  reg [31:0] _RAND_5;
  assign io_out = delays_5; // @[ShiftRegs.scala 24:10:@2814.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delays_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  delays_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delays_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  delays_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  delays_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  delays_5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      delays_0 <= 16'h0;
    end else begin
      delays_0 <= io_in;
    end
    if (reset) begin
      delays_1 <= 16'h0;
    end else begin
      delays_1 <= delays_0;
    end
    if (reset) begin
      delays_2 <= 16'h0;
    end else begin
      delays_2 <= delays_1;
    end
    if (reset) begin
      delays_3 <= 16'h0;
    end else begin
      delays_3 <= delays_2;
    end
    if (reset) begin
      delays_4 <= 16'h0;
    end else begin
      delays_4 <= delays_3;
    end
    if (reset) begin
      delays_5 <= 16'h0;
    end else begin
      delays_5 <= delays_4;
    end
  end
endmodule
module ShiftRegs_6( // @[:@2816.2]
  input         clock, // @[:@2817.4]
  input         reset, // @[:@2818.4]
  input  [15:0] io_in, // @[:@2819.4]
  output [15:0] io_out // @[:@2819.4]
);
  reg [15:0] delays_0; // @[ShiftRegs.scala 15:23:@2829.4]
  reg [31:0] _RAND_0;
  reg [15:0] delays_1; // @[ShiftRegs.scala 15:23:@2829.4]
  reg [31:0] _RAND_1;
  reg [15:0] delays_2; // @[ShiftRegs.scala 15:23:@2829.4]
  reg [31:0] _RAND_2;
  reg [15:0] delays_3; // @[ShiftRegs.scala 15:23:@2829.4]
  reg [31:0] _RAND_3;
  reg [15:0] delays_4; // @[ShiftRegs.scala 15:23:@2829.4]
  reg [31:0] _RAND_4;
  reg [15:0] delays_5; // @[ShiftRegs.scala 15:23:@2829.4]
  reg [31:0] _RAND_5;
  reg [15:0] delays_6; // @[ShiftRegs.scala 15:23:@2829.4]
  reg [31:0] _RAND_6;
  assign io_out = delays_6; // @[ShiftRegs.scala 24:10:@2837.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delays_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  delays_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delays_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  delays_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  delays_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  delays_5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  delays_6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      delays_0 <= 16'h0;
    end else begin
      delays_0 <= io_in;
    end
    if (reset) begin
      delays_1 <= 16'h0;
    end else begin
      delays_1 <= delays_0;
    end
    if (reset) begin
      delays_2 <= 16'h0;
    end else begin
      delays_2 <= delays_1;
    end
    if (reset) begin
      delays_3 <= 16'h0;
    end else begin
      delays_3 <= delays_2;
    end
    if (reset) begin
      delays_4 <= 16'h0;
    end else begin
      delays_4 <= delays_3;
    end
    if (reset) begin
      delays_5 <= 16'h0;
    end else begin
      delays_5 <= delays_4;
    end
    if (reset) begin
      delays_6 <= 16'h0;
    end else begin
      delays_6 <= delays_5;
    end
  end
endmodule
module ShiftRegs_7( // @[:@2839.2]
  input         clock, // @[:@2840.4]
  input         reset, // @[:@2841.4]
  input  [15:0] io_in, // @[:@2842.4]
  output [15:0] io_out // @[:@2842.4]
);
  reg [15:0] delays_0; // @[ShiftRegs.scala 15:23:@2853.4]
  reg [31:0] _RAND_0;
  reg [15:0] delays_1; // @[ShiftRegs.scala 15:23:@2853.4]
  reg [31:0] _RAND_1;
  reg [15:0] delays_2; // @[ShiftRegs.scala 15:23:@2853.4]
  reg [31:0] _RAND_2;
  reg [15:0] delays_3; // @[ShiftRegs.scala 15:23:@2853.4]
  reg [31:0] _RAND_3;
  reg [15:0] delays_4; // @[ShiftRegs.scala 15:23:@2853.4]
  reg [31:0] _RAND_4;
  reg [15:0] delays_5; // @[ShiftRegs.scala 15:23:@2853.4]
  reg [31:0] _RAND_5;
  reg [15:0] delays_6; // @[ShiftRegs.scala 15:23:@2853.4]
  reg [31:0] _RAND_6;
  reg [15:0] delays_7; // @[ShiftRegs.scala 15:23:@2853.4]
  reg [31:0] _RAND_7;
  assign io_out = delays_7; // @[ShiftRegs.scala 24:10:@2862.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delays_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  delays_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delays_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  delays_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  delays_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  delays_5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  delays_6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  delays_7 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      delays_0 <= 16'h0;
    end else begin
      delays_0 <= io_in;
    end
    if (reset) begin
      delays_1 <= 16'h0;
    end else begin
      delays_1 <= delays_0;
    end
    if (reset) begin
      delays_2 <= 16'h0;
    end else begin
      delays_2 <= delays_1;
    end
    if (reset) begin
      delays_3 <= 16'h0;
    end else begin
      delays_3 <= delays_2;
    end
    if (reset) begin
      delays_4 <= 16'h0;
    end else begin
      delays_4 <= delays_3;
    end
    if (reset) begin
      delays_5 <= 16'h0;
    end else begin
      delays_5 <= delays_4;
    end
    if (reset) begin
      delays_6 <= 16'h0;
    end else begin
      delays_6 <= delays_5;
    end
    if (reset) begin
      delays_7 <= 16'h0;
    end else begin
      delays_7 <= delays_6;
    end
  end
endmodule
module ShiftRegs_8( // @[:@2864.2]
  input         clock, // @[:@2865.4]
  input         reset, // @[:@2866.4]
  input  [15:0] io_in, // @[:@2867.4]
  output [15:0] io_out // @[:@2867.4]
);
  reg [15:0] delays_0; // @[ShiftRegs.scala 15:23:@2879.4]
  reg [31:0] _RAND_0;
  reg [15:0] delays_1; // @[ShiftRegs.scala 15:23:@2879.4]
  reg [31:0] _RAND_1;
  reg [15:0] delays_2; // @[ShiftRegs.scala 15:23:@2879.4]
  reg [31:0] _RAND_2;
  reg [15:0] delays_3; // @[ShiftRegs.scala 15:23:@2879.4]
  reg [31:0] _RAND_3;
  reg [15:0] delays_4; // @[ShiftRegs.scala 15:23:@2879.4]
  reg [31:0] _RAND_4;
  reg [15:0] delays_5; // @[ShiftRegs.scala 15:23:@2879.4]
  reg [31:0] _RAND_5;
  reg [15:0] delays_6; // @[ShiftRegs.scala 15:23:@2879.4]
  reg [31:0] _RAND_6;
  reg [15:0] delays_7; // @[ShiftRegs.scala 15:23:@2879.4]
  reg [31:0] _RAND_7;
  reg [15:0] delays_8; // @[ShiftRegs.scala 15:23:@2879.4]
  reg [31:0] _RAND_8;
  assign io_out = delays_8; // @[ShiftRegs.scala 24:10:@2889.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delays_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  delays_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delays_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  delays_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  delays_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  delays_5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  delays_6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  delays_7 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  delays_8 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      delays_0 <= 16'h0;
    end else begin
      delays_0 <= io_in;
    end
    if (reset) begin
      delays_1 <= 16'h0;
    end else begin
      delays_1 <= delays_0;
    end
    if (reset) begin
      delays_2 <= 16'h0;
    end else begin
      delays_2 <= delays_1;
    end
    if (reset) begin
      delays_3 <= 16'h0;
    end else begin
      delays_3 <= delays_2;
    end
    if (reset) begin
      delays_4 <= 16'h0;
    end else begin
      delays_4 <= delays_3;
    end
    if (reset) begin
      delays_5 <= 16'h0;
    end else begin
      delays_5 <= delays_4;
    end
    if (reset) begin
      delays_6 <= 16'h0;
    end else begin
      delays_6 <= delays_5;
    end
    if (reset) begin
      delays_7 <= 16'h0;
    end else begin
      delays_7 <= delays_6;
    end
    if (reset) begin
      delays_8 <= 16'h0;
    end else begin
      delays_8 <= delays_7;
    end
  end
endmodule
module ShiftRegs_9( // @[:@2891.2]
  input         clock, // @[:@2892.4]
  input         reset, // @[:@2893.4]
  input  [15:0] io_in, // @[:@2894.4]
  output [15:0] io_out // @[:@2894.4]
);
  reg [15:0] delays_0; // @[ShiftRegs.scala 15:23:@2907.4]
  reg [31:0] _RAND_0;
  reg [15:0] delays_1; // @[ShiftRegs.scala 15:23:@2907.4]
  reg [31:0] _RAND_1;
  reg [15:0] delays_2; // @[ShiftRegs.scala 15:23:@2907.4]
  reg [31:0] _RAND_2;
  reg [15:0] delays_3; // @[ShiftRegs.scala 15:23:@2907.4]
  reg [31:0] _RAND_3;
  reg [15:0] delays_4; // @[ShiftRegs.scala 15:23:@2907.4]
  reg [31:0] _RAND_4;
  reg [15:0] delays_5; // @[ShiftRegs.scala 15:23:@2907.4]
  reg [31:0] _RAND_5;
  reg [15:0] delays_6; // @[ShiftRegs.scala 15:23:@2907.4]
  reg [31:0] _RAND_6;
  reg [15:0] delays_7; // @[ShiftRegs.scala 15:23:@2907.4]
  reg [31:0] _RAND_7;
  reg [15:0] delays_8; // @[ShiftRegs.scala 15:23:@2907.4]
  reg [31:0] _RAND_8;
  reg [15:0] delays_9; // @[ShiftRegs.scala 15:23:@2907.4]
  reg [31:0] _RAND_9;
  assign io_out = delays_9; // @[ShiftRegs.scala 24:10:@2918.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delays_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  delays_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delays_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  delays_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  delays_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  delays_5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  delays_6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  delays_7 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  delays_8 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  delays_9 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      delays_0 <= 16'h0;
    end else begin
      delays_0 <= io_in;
    end
    if (reset) begin
      delays_1 <= 16'h0;
    end else begin
      delays_1 <= delays_0;
    end
    if (reset) begin
      delays_2 <= 16'h0;
    end else begin
      delays_2 <= delays_1;
    end
    if (reset) begin
      delays_3 <= 16'h0;
    end else begin
      delays_3 <= delays_2;
    end
    if (reset) begin
      delays_4 <= 16'h0;
    end else begin
      delays_4 <= delays_3;
    end
    if (reset) begin
      delays_5 <= 16'h0;
    end else begin
      delays_5 <= delays_4;
    end
    if (reset) begin
      delays_6 <= 16'h0;
    end else begin
      delays_6 <= delays_5;
    end
    if (reset) begin
      delays_7 <= 16'h0;
    end else begin
      delays_7 <= delays_6;
    end
    if (reset) begin
      delays_8 <= 16'h0;
    end else begin
      delays_8 <= delays_7;
    end
    if (reset) begin
      delays_9 <= 16'h0;
    end else begin
      delays_9 <= delays_8;
    end
  end
endmodule
module MMB( // @[:@2920.2]
  input          clock, // @[:@2921.4]
  input          reset, // @[:@2922.4]
  input  [162:0] io_a, // @[:@2923.4]
  input  [162:0] io_bi, // @[:@2923.4]
  output [162:0] io_pout // @[:@2923.4]
);
  wire  PEAlter_clock; // @[MM.scala 16:59:@2925.4]
  wire [162:0] PEAlter_io_a; // @[MM.scala 16:59:@2925.4]
  wire [162:0] PEAlter_io_p; // @[MM.scala 16:59:@2925.4]
  wire [15:0] PEAlter_io_bi; // @[MM.scala 16:59:@2925.4]
  wire [162:0] PEAlter_io_aout; // @[MM.scala 16:59:@2925.4]
  wire [162:0] PEAlter_io_pout; // @[MM.scala 16:59:@2925.4]
  wire  PEAlter_1_clock; // @[MM.scala 16:59:@2928.4]
  wire [162:0] PEAlter_1_io_a; // @[MM.scala 16:59:@2928.4]
  wire [162:0] PEAlter_1_io_p; // @[MM.scala 16:59:@2928.4]
  wire [15:0] PEAlter_1_io_bi; // @[MM.scala 16:59:@2928.4]
  wire [162:0] PEAlter_1_io_aout; // @[MM.scala 16:59:@2928.4]
  wire [162:0] PEAlter_1_io_pout; // @[MM.scala 16:59:@2928.4]
  wire  PEAlter_2_clock; // @[MM.scala 16:59:@2931.4]
  wire [162:0] PEAlter_2_io_a; // @[MM.scala 16:59:@2931.4]
  wire [162:0] PEAlter_2_io_p; // @[MM.scala 16:59:@2931.4]
  wire [15:0] PEAlter_2_io_bi; // @[MM.scala 16:59:@2931.4]
  wire [162:0] PEAlter_2_io_aout; // @[MM.scala 16:59:@2931.4]
  wire [162:0] PEAlter_2_io_pout; // @[MM.scala 16:59:@2931.4]
  wire  PEAlter_3_clock; // @[MM.scala 16:59:@2934.4]
  wire [162:0] PEAlter_3_io_a; // @[MM.scala 16:59:@2934.4]
  wire [162:0] PEAlter_3_io_p; // @[MM.scala 16:59:@2934.4]
  wire [15:0] PEAlter_3_io_bi; // @[MM.scala 16:59:@2934.4]
  wire [162:0] PEAlter_3_io_aout; // @[MM.scala 16:59:@2934.4]
  wire [162:0] PEAlter_3_io_pout; // @[MM.scala 16:59:@2934.4]
  wire  PEAlter_4_clock; // @[MM.scala 16:59:@2937.4]
  wire [162:0] PEAlter_4_io_a; // @[MM.scala 16:59:@2937.4]
  wire [162:0] PEAlter_4_io_p; // @[MM.scala 16:59:@2937.4]
  wire [15:0] PEAlter_4_io_bi; // @[MM.scala 16:59:@2937.4]
  wire [162:0] PEAlter_4_io_aout; // @[MM.scala 16:59:@2937.4]
  wire [162:0] PEAlter_4_io_pout; // @[MM.scala 16:59:@2937.4]
  wire  PEAlter_5_clock; // @[MM.scala 16:59:@2940.4]
  wire [162:0] PEAlter_5_io_a; // @[MM.scala 16:59:@2940.4]
  wire [162:0] PEAlter_5_io_p; // @[MM.scala 16:59:@2940.4]
  wire [15:0] PEAlter_5_io_bi; // @[MM.scala 16:59:@2940.4]
  wire [162:0] PEAlter_5_io_aout; // @[MM.scala 16:59:@2940.4]
  wire [162:0] PEAlter_5_io_pout; // @[MM.scala 16:59:@2940.4]
  wire  PEAlter_6_clock; // @[MM.scala 16:59:@2943.4]
  wire [162:0] PEAlter_6_io_a; // @[MM.scala 16:59:@2943.4]
  wire [162:0] PEAlter_6_io_p; // @[MM.scala 16:59:@2943.4]
  wire [15:0] PEAlter_6_io_bi; // @[MM.scala 16:59:@2943.4]
  wire [162:0] PEAlter_6_io_aout; // @[MM.scala 16:59:@2943.4]
  wire [162:0] PEAlter_6_io_pout; // @[MM.scala 16:59:@2943.4]
  wire  PEAlter_7_clock; // @[MM.scala 16:59:@2946.4]
  wire [162:0] PEAlter_7_io_a; // @[MM.scala 16:59:@2946.4]
  wire [162:0] PEAlter_7_io_p; // @[MM.scala 16:59:@2946.4]
  wire [15:0] PEAlter_7_io_bi; // @[MM.scala 16:59:@2946.4]
  wire [162:0] PEAlter_7_io_aout; // @[MM.scala 16:59:@2946.4]
  wire [162:0] PEAlter_7_io_pout; // @[MM.scala 16:59:@2946.4]
  wire  PEAlter_8_clock; // @[MM.scala 16:59:@2949.4]
  wire [162:0] PEAlter_8_io_a; // @[MM.scala 16:59:@2949.4]
  wire [162:0] PEAlter_8_io_p; // @[MM.scala 16:59:@2949.4]
  wire [15:0] PEAlter_8_io_bi; // @[MM.scala 16:59:@2949.4]
  wire [162:0] PEAlter_8_io_aout; // @[MM.scala 16:59:@2949.4]
  wire [162:0] PEAlter_8_io_pout; // @[MM.scala 16:59:@2949.4]
  wire  PEAlter_9_clock; // @[MM.scala 16:59:@2952.4]
  wire [162:0] PEAlter_9_io_a; // @[MM.scala 16:59:@2952.4]
  wire [162:0] PEAlter_9_io_p; // @[MM.scala 16:59:@2952.4]
  wire [15:0] PEAlter_9_io_bi; // @[MM.scala 16:59:@2952.4]
  wire [162:0] PEAlter_9_io_aout; // @[MM.scala 16:59:@2952.4]
  wire [162:0] PEAlter_9_io_pout; // @[MM.scala 16:59:@2952.4]
  wire  PEAlter_10_clock; // @[MM.scala 16:59:@2955.4]
  wire [162:0] PEAlter_10_io_a; // @[MM.scala 16:59:@2955.4]
  wire [162:0] PEAlter_10_io_p; // @[MM.scala 16:59:@2955.4]
  wire [15:0] PEAlter_10_io_bi; // @[MM.scala 16:59:@2955.4]
  wire [162:0] PEAlter_10_io_aout; // @[MM.scala 16:59:@2955.4]
  wire [162:0] PEAlter_10_io_pout; // @[MM.scala 16:59:@2955.4]
  wire  ShiftRegs_clock; // @[ShiftRegs.scala 30:22:@3022.4]
  wire  ShiftRegs_reset; // @[ShiftRegs.scala 30:22:@3022.4]
  wire [15:0] ShiftRegs_io_in; // @[ShiftRegs.scala 30:22:@3022.4]
  wire [15:0] ShiftRegs_io_out; // @[ShiftRegs.scala 30:22:@3022.4]
  wire  ShiftRegs_1_clock; // @[ShiftRegs.scala 30:22:@3030.4]
  wire  ShiftRegs_1_reset; // @[ShiftRegs.scala 30:22:@3030.4]
  wire [15:0] ShiftRegs_1_io_in; // @[ShiftRegs.scala 30:22:@3030.4]
  wire [15:0] ShiftRegs_1_io_out; // @[ShiftRegs.scala 30:22:@3030.4]
  wire  ShiftRegs_2_clock; // @[ShiftRegs.scala 30:22:@3038.4]
  wire  ShiftRegs_2_reset; // @[ShiftRegs.scala 30:22:@3038.4]
  wire [15:0] ShiftRegs_2_io_in; // @[ShiftRegs.scala 30:22:@3038.4]
  wire [15:0] ShiftRegs_2_io_out; // @[ShiftRegs.scala 30:22:@3038.4]
  wire  ShiftRegs_3_clock; // @[ShiftRegs.scala 30:22:@3046.4]
  wire  ShiftRegs_3_reset; // @[ShiftRegs.scala 30:22:@3046.4]
  wire [15:0] ShiftRegs_3_io_in; // @[ShiftRegs.scala 30:22:@3046.4]
  wire [15:0] ShiftRegs_3_io_out; // @[ShiftRegs.scala 30:22:@3046.4]
  wire  ShiftRegs_4_clock; // @[ShiftRegs.scala 30:22:@3054.4]
  wire  ShiftRegs_4_reset; // @[ShiftRegs.scala 30:22:@3054.4]
  wire [15:0] ShiftRegs_4_io_in; // @[ShiftRegs.scala 30:22:@3054.4]
  wire [15:0] ShiftRegs_4_io_out; // @[ShiftRegs.scala 30:22:@3054.4]
  wire  ShiftRegs_5_clock; // @[ShiftRegs.scala 30:22:@3062.4]
  wire  ShiftRegs_5_reset; // @[ShiftRegs.scala 30:22:@3062.4]
  wire [15:0] ShiftRegs_5_io_in; // @[ShiftRegs.scala 30:22:@3062.4]
  wire [15:0] ShiftRegs_5_io_out; // @[ShiftRegs.scala 30:22:@3062.4]
  wire  ShiftRegs_6_clock; // @[ShiftRegs.scala 30:22:@3070.4]
  wire  ShiftRegs_6_reset; // @[ShiftRegs.scala 30:22:@3070.4]
  wire [15:0] ShiftRegs_6_io_in; // @[ShiftRegs.scala 30:22:@3070.4]
  wire [15:0] ShiftRegs_6_io_out; // @[ShiftRegs.scala 30:22:@3070.4]
  wire  ShiftRegs_7_clock; // @[ShiftRegs.scala 30:22:@3078.4]
  wire  ShiftRegs_7_reset; // @[ShiftRegs.scala 30:22:@3078.4]
  wire [15:0] ShiftRegs_7_io_in; // @[ShiftRegs.scala 30:22:@3078.4]
  wire [15:0] ShiftRegs_7_io_out; // @[ShiftRegs.scala 30:22:@3078.4]
  wire  ShiftRegs_8_clock; // @[ShiftRegs.scala 30:22:@3086.4]
  wire  ShiftRegs_8_reset; // @[ShiftRegs.scala 30:22:@3086.4]
  wire [15:0] ShiftRegs_8_io_in; // @[ShiftRegs.scala 30:22:@3086.4]
  wire [15:0] ShiftRegs_8_io_out; // @[ShiftRegs.scala 30:22:@3086.4]
  wire  ShiftRegs_9_clock; // @[ShiftRegs.scala 30:22:@3094.4]
  wire  ShiftRegs_9_reset; // @[ShiftRegs.scala 30:22:@3094.4]
  wire [15:0] ShiftRegs_9_io_in; // @[ShiftRegs.scala 30:22:@3094.4]
  wire [15:0] ShiftRegs_9_io_out; // @[ShiftRegs.scala 30:22:@3094.4]
  wire [2:0] _T_215; // @[MM.scala 22:52:@3016.4]
  PEAlter PEAlter ( // @[MM.scala 16:59:@2925.4]
    .clock(PEAlter_clock),
    .io_a(PEAlter_io_a),
    .io_p(PEAlter_io_p),
    .io_bi(PEAlter_io_bi),
    .io_aout(PEAlter_io_aout),
    .io_pout(PEAlter_io_pout)
  );
  PEAlter PEAlter_1 ( // @[MM.scala 16:59:@2928.4]
    .clock(PEAlter_1_clock),
    .io_a(PEAlter_1_io_a),
    .io_p(PEAlter_1_io_p),
    .io_bi(PEAlter_1_io_bi),
    .io_aout(PEAlter_1_io_aout),
    .io_pout(PEAlter_1_io_pout)
  );
  PEAlter PEAlter_2 ( // @[MM.scala 16:59:@2931.4]
    .clock(PEAlter_2_clock),
    .io_a(PEAlter_2_io_a),
    .io_p(PEAlter_2_io_p),
    .io_bi(PEAlter_2_io_bi),
    .io_aout(PEAlter_2_io_aout),
    .io_pout(PEAlter_2_io_pout)
  );
  PEAlter PEAlter_3 ( // @[MM.scala 16:59:@2934.4]
    .clock(PEAlter_3_clock),
    .io_a(PEAlter_3_io_a),
    .io_p(PEAlter_3_io_p),
    .io_bi(PEAlter_3_io_bi),
    .io_aout(PEAlter_3_io_aout),
    .io_pout(PEAlter_3_io_pout)
  );
  PEAlter PEAlter_4 ( // @[MM.scala 16:59:@2937.4]
    .clock(PEAlter_4_clock),
    .io_a(PEAlter_4_io_a),
    .io_p(PEAlter_4_io_p),
    .io_bi(PEAlter_4_io_bi),
    .io_aout(PEAlter_4_io_aout),
    .io_pout(PEAlter_4_io_pout)
  );
  PEAlter PEAlter_5 ( // @[MM.scala 16:59:@2940.4]
    .clock(PEAlter_5_clock),
    .io_a(PEAlter_5_io_a),
    .io_p(PEAlter_5_io_p),
    .io_bi(PEAlter_5_io_bi),
    .io_aout(PEAlter_5_io_aout),
    .io_pout(PEAlter_5_io_pout)
  );
  PEAlter PEAlter_6 ( // @[MM.scala 16:59:@2943.4]
    .clock(PEAlter_6_clock),
    .io_a(PEAlter_6_io_a),
    .io_p(PEAlter_6_io_p),
    .io_bi(PEAlter_6_io_bi),
    .io_aout(PEAlter_6_io_aout),
    .io_pout(PEAlter_6_io_pout)
  );
  PEAlter PEAlter_7 ( // @[MM.scala 16:59:@2946.4]
    .clock(PEAlter_7_clock),
    .io_a(PEAlter_7_io_a),
    .io_p(PEAlter_7_io_p),
    .io_bi(PEAlter_7_io_bi),
    .io_aout(PEAlter_7_io_aout),
    .io_pout(PEAlter_7_io_pout)
  );
  PEAlter PEAlter_8 ( // @[MM.scala 16:59:@2949.4]
    .clock(PEAlter_8_clock),
    .io_a(PEAlter_8_io_a),
    .io_p(PEAlter_8_io_p),
    .io_bi(PEAlter_8_io_bi),
    .io_aout(PEAlter_8_io_aout),
    .io_pout(PEAlter_8_io_pout)
  );
  PEAlter PEAlter_9 ( // @[MM.scala 16:59:@2952.4]
    .clock(PEAlter_9_clock),
    .io_a(PEAlter_9_io_a),
    .io_p(PEAlter_9_io_p),
    .io_bi(PEAlter_9_io_bi),
    .io_aout(PEAlter_9_io_aout),
    .io_pout(PEAlter_9_io_pout)
  );
  PEAlter PEAlter_10 ( // @[MM.scala 16:59:@2955.4]
    .clock(PEAlter_10_clock),
    .io_a(PEAlter_10_io_a),
    .io_p(PEAlter_10_io_p),
    .io_bi(PEAlter_10_io_bi),
    .io_aout(PEAlter_10_io_aout),
    .io_pout(PEAlter_10_io_pout)
  );
  ShiftRegs ShiftRegs ( // @[ShiftRegs.scala 30:22:@3022.4]
    .clock(ShiftRegs_clock),
    .reset(ShiftRegs_reset),
    .io_in(ShiftRegs_io_in),
    .io_out(ShiftRegs_io_out)
  );
  ShiftRegs_1 ShiftRegs_1 ( // @[ShiftRegs.scala 30:22:@3030.4]
    .clock(ShiftRegs_1_clock),
    .reset(ShiftRegs_1_reset),
    .io_in(ShiftRegs_1_io_in),
    .io_out(ShiftRegs_1_io_out)
  );
  ShiftRegs_2 ShiftRegs_2 ( // @[ShiftRegs.scala 30:22:@3038.4]
    .clock(ShiftRegs_2_clock),
    .reset(ShiftRegs_2_reset),
    .io_in(ShiftRegs_2_io_in),
    .io_out(ShiftRegs_2_io_out)
  );
  ShiftRegs_3 ShiftRegs_3 ( // @[ShiftRegs.scala 30:22:@3046.4]
    .clock(ShiftRegs_3_clock),
    .reset(ShiftRegs_3_reset),
    .io_in(ShiftRegs_3_io_in),
    .io_out(ShiftRegs_3_io_out)
  );
  ShiftRegs_4 ShiftRegs_4 ( // @[ShiftRegs.scala 30:22:@3054.4]
    .clock(ShiftRegs_4_clock),
    .reset(ShiftRegs_4_reset),
    .io_in(ShiftRegs_4_io_in),
    .io_out(ShiftRegs_4_io_out)
  );
  ShiftRegs_5 ShiftRegs_5 ( // @[ShiftRegs.scala 30:22:@3062.4]
    .clock(ShiftRegs_5_clock),
    .reset(ShiftRegs_5_reset),
    .io_in(ShiftRegs_5_io_in),
    .io_out(ShiftRegs_5_io_out)
  );
  ShiftRegs_6 ShiftRegs_6 ( // @[ShiftRegs.scala 30:22:@3070.4]
    .clock(ShiftRegs_6_clock),
    .reset(ShiftRegs_6_reset),
    .io_in(ShiftRegs_6_io_in),
    .io_out(ShiftRegs_6_io_out)
  );
  ShiftRegs_7 ShiftRegs_7 ( // @[ShiftRegs.scala 30:22:@3078.4]
    .clock(ShiftRegs_7_clock),
    .reset(ShiftRegs_7_reset),
    .io_in(ShiftRegs_7_io_in),
    .io_out(ShiftRegs_7_io_out)
  );
  ShiftRegs_8 ShiftRegs_8 ( // @[ShiftRegs.scala 30:22:@3086.4]
    .clock(ShiftRegs_8_clock),
    .reset(ShiftRegs_8_reset),
    .io_in(ShiftRegs_8_io_in),
    .io_out(ShiftRegs_8_io_out)
  );
  ShiftRegs_9 ShiftRegs_9 ( // @[ShiftRegs.scala 30:22:@3094.4]
    .clock(ShiftRegs_9_clock),
    .reset(ShiftRegs_9_reset),
    .io_in(ShiftRegs_9_io_in),
    .io_out(ShiftRegs_9_io_out)
  );
  assign _T_215 = io_bi[162:160]; // @[MM.scala 22:52:@3016.4]
  assign io_pout = PEAlter_10_io_pout; // @[MM.scala 31:13:@3099.4]
  assign PEAlter_clock = clock; // @[:@2926.4]
  assign PEAlter_io_a = io_a; // @[MM.scala 16:22:@2963.4]
  assign PEAlter_io_p = 163'h0; // @[MM.scala 16:22:@2962.4]
  assign PEAlter_io_bi = {13'h0,_T_215}; // @[MM.scala 16:22:@2961.4]
  assign PEAlter_1_clock = clock; // @[:@2929.4]
  assign PEAlter_1_io_a = PEAlter_io_aout; // @[MM.scala 16:22:@2968.4]
  assign PEAlter_1_io_p = PEAlter_io_pout; // @[MM.scala 16:22:@2967.4]
  assign PEAlter_1_io_bi = ShiftRegs_io_out; // @[MM.scala 16:22:@2966.4]
  assign PEAlter_2_clock = clock; // @[:@2932.4]
  assign PEAlter_2_io_a = PEAlter_1_io_aout; // @[MM.scala 16:22:@2973.4]
  assign PEAlter_2_io_p = PEAlter_1_io_pout; // @[MM.scala 16:22:@2972.4]
  assign PEAlter_2_io_bi = ShiftRegs_1_io_out; // @[MM.scala 16:22:@2971.4]
  assign PEAlter_3_clock = clock; // @[:@2935.4]
  assign PEAlter_3_io_a = PEAlter_2_io_aout; // @[MM.scala 16:22:@2978.4]
  assign PEAlter_3_io_p = PEAlter_2_io_pout; // @[MM.scala 16:22:@2977.4]
  assign PEAlter_3_io_bi = ShiftRegs_2_io_out; // @[MM.scala 16:22:@2976.4]
  assign PEAlter_4_clock = clock; // @[:@2938.4]
  assign PEAlter_4_io_a = PEAlter_3_io_aout; // @[MM.scala 16:22:@2983.4]
  assign PEAlter_4_io_p = PEAlter_3_io_pout; // @[MM.scala 16:22:@2982.4]
  assign PEAlter_4_io_bi = ShiftRegs_3_io_out; // @[MM.scala 16:22:@2981.4]
  assign PEAlter_5_clock = clock; // @[:@2941.4]
  assign PEAlter_5_io_a = PEAlter_4_io_aout; // @[MM.scala 16:22:@2988.4]
  assign PEAlter_5_io_p = PEAlter_4_io_pout; // @[MM.scala 16:22:@2987.4]
  assign PEAlter_5_io_bi = ShiftRegs_4_io_out; // @[MM.scala 16:22:@2986.4]
  assign PEAlter_6_clock = clock; // @[:@2944.4]
  assign PEAlter_6_io_a = PEAlter_5_io_aout; // @[MM.scala 16:22:@2993.4]
  assign PEAlter_6_io_p = PEAlter_5_io_pout; // @[MM.scala 16:22:@2992.4]
  assign PEAlter_6_io_bi = ShiftRegs_5_io_out; // @[MM.scala 16:22:@2991.4]
  assign PEAlter_7_clock = clock; // @[:@2947.4]
  assign PEAlter_7_io_a = PEAlter_6_io_aout; // @[MM.scala 16:22:@2998.4]
  assign PEAlter_7_io_p = PEAlter_6_io_pout; // @[MM.scala 16:22:@2997.4]
  assign PEAlter_7_io_bi = ShiftRegs_6_io_out; // @[MM.scala 16:22:@2996.4]
  assign PEAlter_8_clock = clock; // @[:@2950.4]
  assign PEAlter_8_io_a = PEAlter_7_io_aout; // @[MM.scala 16:22:@3003.4]
  assign PEAlter_8_io_p = PEAlter_7_io_pout; // @[MM.scala 16:22:@3002.4]
  assign PEAlter_8_io_bi = ShiftRegs_7_io_out; // @[MM.scala 16:22:@3001.4]
  assign PEAlter_9_clock = clock; // @[:@2953.4]
  assign PEAlter_9_io_a = PEAlter_8_io_aout; // @[MM.scala 16:22:@3008.4]
  assign PEAlter_9_io_p = PEAlter_8_io_pout; // @[MM.scala 16:22:@3007.4]
  assign PEAlter_9_io_bi = ShiftRegs_8_io_out; // @[MM.scala 16:22:@3006.4]
  assign PEAlter_10_clock = clock; // @[:@2956.4]
  assign PEAlter_10_io_a = PEAlter_9_io_aout; // @[MM.scala 16:22:@3013.4]
  assign PEAlter_10_io_p = PEAlter_9_io_pout; // @[MM.scala 16:22:@3012.4]
  assign PEAlter_10_io_bi = ShiftRegs_9_io_out; // @[MM.scala 16:22:@3011.4]
  assign ShiftRegs_clock = clock; // @[:@3023.4]
  assign ShiftRegs_reset = reset; // @[:@3024.4]
  assign ShiftRegs_io_in = io_bi[159:144]; // @[ShiftRegs.scala 31:16:@3025.4]
  assign ShiftRegs_1_clock = clock; // @[:@3031.4]
  assign ShiftRegs_1_reset = reset; // @[:@3032.4]
  assign ShiftRegs_1_io_in = io_bi[143:128]; // @[ShiftRegs.scala 31:16:@3033.4]
  assign ShiftRegs_2_clock = clock; // @[:@3039.4]
  assign ShiftRegs_2_reset = reset; // @[:@3040.4]
  assign ShiftRegs_2_io_in = io_bi[127:112]; // @[ShiftRegs.scala 31:16:@3041.4]
  assign ShiftRegs_3_clock = clock; // @[:@3047.4]
  assign ShiftRegs_3_reset = reset; // @[:@3048.4]
  assign ShiftRegs_3_io_in = io_bi[111:96]; // @[ShiftRegs.scala 31:16:@3049.4]
  assign ShiftRegs_4_clock = clock; // @[:@3055.4]
  assign ShiftRegs_4_reset = reset; // @[:@3056.4]
  assign ShiftRegs_4_io_in = io_bi[95:80]; // @[ShiftRegs.scala 31:16:@3057.4]
  assign ShiftRegs_5_clock = clock; // @[:@3063.4]
  assign ShiftRegs_5_reset = reset; // @[:@3064.4]
  assign ShiftRegs_5_io_in = io_bi[79:64]; // @[ShiftRegs.scala 31:16:@3065.4]
  assign ShiftRegs_6_clock = clock; // @[:@3071.4]
  assign ShiftRegs_6_reset = reset; // @[:@3072.4]
  assign ShiftRegs_6_io_in = io_bi[63:48]; // @[ShiftRegs.scala 31:16:@3073.4]
  assign ShiftRegs_7_clock = clock; // @[:@3079.4]
  assign ShiftRegs_7_reset = reset; // @[:@3080.4]
  assign ShiftRegs_7_io_in = io_bi[47:32]; // @[ShiftRegs.scala 31:16:@3081.4]
  assign ShiftRegs_8_clock = clock; // @[:@3087.4]
  assign ShiftRegs_8_reset = reset; // @[:@3088.4]
  assign ShiftRegs_8_io_in = io_bi[31:16]; // @[ShiftRegs.scala 31:16:@3089.4]
  assign ShiftRegs_9_clock = clock; // @[:@3095.4]
  assign ShiftRegs_9_reset = reset; // @[:@3096.4]
  assign ShiftRegs_9_io_in = io_bi[15:0]; // @[ShiftRegs.scala 31:16:@3097.4]
endmodule
