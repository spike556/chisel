module FMul( // @[:@3.2]
  input  [162:0] io_a, // @[:@6.4]
  input  [31:0]  io_b, // @[:@6.4]
  output [193:0] io_pout // @[:@6.4]
);
  wire  _T_148; // @[PEAlter.scala 19:15:@108.4]
  wire [163:0] _GEN_32; // @[PEAlter.scala 20:34:@111.6]
  wire [163:0] _T_152; // @[PEAlter.scala 20:34:@111.6]
  wire [193:0] _T_153; // @[PEAlter.scala 20:26:@112.6]
  wire [193:0] tmp_1; // @[PEAlter.scala 19:28:@110.4]
  wire  _T_154; // @[PEAlter.scala 19:15:@118.4]
  wire [163:0] _T_158; // @[PEAlter.scala 20:34:@121.6]
  wire [193:0] _GEN_34; // @[PEAlter.scala 20:26:@122.6]
  wire [193:0] _T_159; // @[PEAlter.scala 20:26:@122.6]
  wire [193:0] tmp_2; // @[PEAlter.scala 19:28:@120.4]
  wire  _T_160; // @[PEAlter.scala 19:15:@128.4]
  wire [165:0] _GEN_35; // @[PEAlter.scala 20:34:@131.6]
  wire [165:0] _T_164; // @[PEAlter.scala 20:34:@131.6]
  wire [193:0] _GEN_36; // @[PEAlter.scala 20:26:@132.6]
  wire [193:0] _T_165; // @[PEAlter.scala 20:26:@132.6]
  wire [193:0] tmp_3; // @[PEAlter.scala 19:28:@130.4]
  wire  _T_166; // @[PEAlter.scala 19:15:@138.4]
  wire [165:0] _T_170; // @[PEAlter.scala 20:34:@141.6]
  wire [193:0] _GEN_38; // @[PEAlter.scala 20:26:@142.6]
  wire [193:0] _T_171; // @[PEAlter.scala 20:26:@142.6]
  wire [193:0] tmp_4; // @[PEAlter.scala 19:28:@140.4]
  wire  _T_172; // @[PEAlter.scala 19:15:@148.4]
  wire [169:0] _GEN_39; // @[PEAlter.scala 20:34:@151.6]
  wire [169:0] _T_176; // @[PEAlter.scala 20:34:@151.6]
  wire [193:0] _GEN_40; // @[PEAlter.scala 20:26:@152.6]
  wire [193:0] _T_177; // @[PEAlter.scala 20:26:@152.6]
  wire [193:0] tmp_5; // @[PEAlter.scala 19:28:@150.4]
  wire  _T_178; // @[PEAlter.scala 19:15:@158.4]
  wire [169:0] _T_182; // @[PEAlter.scala 20:34:@161.6]
  wire [193:0] _GEN_42; // @[PEAlter.scala 20:26:@162.6]
  wire [193:0] _T_183; // @[PEAlter.scala 20:26:@162.6]
  wire [193:0] tmp_6; // @[PEAlter.scala 19:28:@160.4]
  wire  _T_184; // @[PEAlter.scala 19:15:@168.4]
  wire [169:0] _T_188; // @[PEAlter.scala 20:34:@171.6]
  wire [193:0] _GEN_44; // @[PEAlter.scala 20:26:@172.6]
  wire [193:0] _T_189; // @[PEAlter.scala 20:26:@172.6]
  wire [193:0] tmp_7; // @[PEAlter.scala 19:28:@170.4]
  wire  _T_190; // @[PEAlter.scala 19:15:@178.4]
  wire [169:0] _T_194; // @[PEAlter.scala 20:34:@181.6]
  wire [193:0] _GEN_46; // @[PEAlter.scala 20:26:@182.6]
  wire [193:0] _T_195; // @[PEAlter.scala 20:26:@182.6]
  wire [193:0] tmp_8; // @[PEAlter.scala 19:28:@180.4]
  wire  _T_196; // @[PEAlter.scala 19:15:@188.4]
  wire [177:0] _GEN_47; // @[PEAlter.scala 20:34:@191.6]
  wire [177:0] _T_200; // @[PEAlter.scala 20:34:@191.6]
  wire [193:0] _GEN_48; // @[PEAlter.scala 20:26:@192.6]
  wire [193:0] _T_201; // @[PEAlter.scala 20:26:@192.6]
  wire [193:0] tmp_9; // @[PEAlter.scala 19:28:@190.4]
  wire  _T_202; // @[PEAlter.scala 19:15:@198.4]
  wire [177:0] _T_206; // @[PEAlter.scala 20:34:@201.6]
  wire [193:0] _GEN_50; // @[PEAlter.scala 20:26:@202.6]
  wire [193:0] _T_207; // @[PEAlter.scala 20:26:@202.6]
  wire [193:0] tmp_10; // @[PEAlter.scala 19:28:@200.4]
  wire  _T_208; // @[PEAlter.scala 19:15:@208.4]
  wire [177:0] _T_212; // @[PEAlter.scala 20:34:@211.6]
  wire [193:0] _GEN_52; // @[PEAlter.scala 20:26:@212.6]
  wire [193:0] _T_213; // @[PEAlter.scala 20:26:@212.6]
  wire [193:0] tmp_11; // @[PEAlter.scala 19:28:@210.4]
  wire  _T_214; // @[PEAlter.scala 19:15:@218.4]
  wire [177:0] _T_218; // @[PEAlter.scala 20:34:@221.6]
  wire [193:0] _GEN_54; // @[PEAlter.scala 20:26:@222.6]
  wire [193:0] _T_219; // @[PEAlter.scala 20:26:@222.6]
  wire [193:0] tmp_12; // @[PEAlter.scala 19:28:@220.4]
  wire  _T_220; // @[PEAlter.scala 19:15:@228.4]
  wire [177:0] _T_224; // @[PEAlter.scala 20:34:@231.6]
  wire [193:0] _GEN_56; // @[PEAlter.scala 20:26:@232.6]
  wire [193:0] _T_225; // @[PEAlter.scala 20:26:@232.6]
  wire [193:0] tmp_13; // @[PEAlter.scala 19:28:@230.4]
  wire  _T_226; // @[PEAlter.scala 19:15:@238.4]
  wire [177:0] _T_230; // @[PEAlter.scala 20:34:@241.6]
  wire [193:0] _GEN_58; // @[PEAlter.scala 20:26:@242.6]
  wire [193:0] _T_231; // @[PEAlter.scala 20:26:@242.6]
  wire [193:0] tmp_14; // @[PEAlter.scala 19:28:@240.4]
  wire  _T_232; // @[PEAlter.scala 19:15:@248.4]
  wire [177:0] _T_236; // @[PEAlter.scala 20:34:@251.6]
  wire [193:0] _GEN_60; // @[PEAlter.scala 20:26:@252.6]
  wire [193:0] _T_237; // @[PEAlter.scala 20:26:@252.6]
  wire [193:0] tmp_15; // @[PEAlter.scala 19:28:@250.4]
  wire  _T_238; // @[PEAlter.scala 19:15:@258.4]
  wire [177:0] _T_242; // @[PEAlter.scala 20:34:@261.6]
  wire [193:0] _GEN_62; // @[PEAlter.scala 20:26:@262.6]
  wire [193:0] _T_243; // @[PEAlter.scala 20:26:@262.6]
  wire [193:0] tmp_16; // @[PEAlter.scala 19:28:@260.4]
  wire  _T_244; // @[PEAlter.scala 19:15:@268.4]
  wire [193:0] _GEN_63; // @[PEAlter.scala 20:34:@271.6]
  wire [193:0] _T_248; // @[PEAlter.scala 20:34:@271.6]
  wire [193:0] _T_249; // @[PEAlter.scala 20:26:@272.6]
  wire [193:0] tmp_17; // @[PEAlter.scala 19:28:@270.4]
  wire  _T_250; // @[PEAlter.scala 19:15:@278.4]
  wire [193:0] _T_254; // @[PEAlter.scala 20:34:@281.6]
  wire [193:0] _T_255; // @[PEAlter.scala 20:26:@282.6]
  wire [193:0] tmp_18; // @[PEAlter.scala 19:28:@280.4]
  wire  _T_256; // @[PEAlter.scala 19:15:@288.4]
  wire [193:0] _T_260; // @[PEAlter.scala 20:34:@291.6]
  wire [193:0] _T_261; // @[PEAlter.scala 20:26:@292.6]
  wire [193:0] tmp_19; // @[PEAlter.scala 19:28:@290.4]
  wire  _T_262; // @[PEAlter.scala 19:15:@298.4]
  wire [193:0] _T_266; // @[PEAlter.scala 20:34:@301.6]
  wire [193:0] _T_267; // @[PEAlter.scala 20:26:@302.6]
  wire [193:0] tmp_20; // @[PEAlter.scala 19:28:@300.4]
  wire  _T_268; // @[PEAlter.scala 19:15:@308.4]
  wire [193:0] _T_272; // @[PEAlter.scala 20:34:@311.6]
  wire [193:0] _T_273; // @[PEAlter.scala 20:26:@312.6]
  wire [193:0] tmp_21; // @[PEAlter.scala 19:28:@310.4]
  wire  _T_274; // @[PEAlter.scala 19:15:@318.4]
  wire [193:0] _T_278; // @[PEAlter.scala 20:34:@321.6]
  wire [193:0] _T_279; // @[PEAlter.scala 20:26:@322.6]
  wire [193:0] tmp_22; // @[PEAlter.scala 19:28:@320.4]
  wire  _T_280; // @[PEAlter.scala 19:15:@328.4]
  wire [193:0] _T_284; // @[PEAlter.scala 20:34:@331.6]
  wire [193:0] _T_285; // @[PEAlter.scala 20:26:@332.6]
  wire [193:0] tmp_23; // @[PEAlter.scala 19:28:@330.4]
  wire  _T_286; // @[PEAlter.scala 19:15:@338.4]
  wire [193:0] _T_290; // @[PEAlter.scala 20:34:@341.6]
  wire [193:0] _T_291; // @[PEAlter.scala 20:26:@342.6]
  wire [193:0] tmp_24; // @[PEAlter.scala 19:28:@340.4]
  wire  _T_292; // @[PEAlter.scala 19:15:@348.4]
  wire [193:0] _T_296; // @[PEAlter.scala 20:34:@351.6]
  wire [193:0] _T_297; // @[PEAlter.scala 20:26:@352.6]
  wire [193:0] tmp_25; // @[PEAlter.scala 19:28:@350.4]
  wire  _T_298; // @[PEAlter.scala 19:15:@358.4]
  wire [193:0] _T_302; // @[PEAlter.scala 20:34:@361.6]
  wire [193:0] _T_303; // @[PEAlter.scala 20:26:@362.6]
  wire [193:0] tmp_26; // @[PEAlter.scala 19:28:@360.4]
  wire  _T_304; // @[PEAlter.scala 19:15:@368.4]
  wire [193:0] _T_308; // @[PEAlter.scala 20:34:@371.6]
  wire [193:0] _T_309; // @[PEAlter.scala 20:26:@372.6]
  wire [193:0] tmp_27; // @[PEAlter.scala 19:28:@370.4]
  wire  _T_310; // @[PEAlter.scala 19:15:@378.4]
  wire [193:0] _T_314; // @[PEAlter.scala 20:34:@381.6]
  wire [193:0] _T_315; // @[PEAlter.scala 20:26:@382.6]
  wire [193:0] tmp_28; // @[PEAlter.scala 19:28:@380.4]
  wire  _T_316; // @[PEAlter.scala 19:15:@388.4]
  wire [193:0] _T_320; // @[PEAlter.scala 20:34:@391.6]
  wire [193:0] _T_321; // @[PEAlter.scala 20:26:@392.6]
  wire [193:0] tmp_29; // @[PEAlter.scala 19:28:@390.4]
  wire  _T_322; // @[PEAlter.scala 19:15:@398.4]
  wire [193:0] _T_326; // @[PEAlter.scala 20:34:@401.6]
  wire [193:0] _T_327; // @[PEAlter.scala 20:26:@402.6]
  wire [193:0] tmp_30; // @[PEAlter.scala 19:28:@400.4]
  wire  _T_328; // @[PEAlter.scala 19:15:@408.4]
  wire [193:0] _T_332; // @[PEAlter.scala 20:34:@411.6]
  wire [193:0] _T_333; // @[PEAlter.scala 20:26:@412.6]
  wire [193:0] tmp_31; // @[PEAlter.scala 19:28:@410.4]
  wire  _T_334; // @[PEAlter.scala 19:15:@418.4]
  wire [193:0] _T_338; // @[PEAlter.scala 20:34:@421.6]
  wire [193:0] _T_339; // @[PEAlter.scala 20:26:@422.6]
  assign _T_148 = io_b[0]; // @[PEAlter.scala 19:15:@108.4]
  assign _GEN_32 = {{1'd0}, io_a}; // @[PEAlter.scala 20:34:@111.6]
  assign _T_152 = _GEN_32 << 1'h0; // @[PEAlter.scala 20:34:@111.6]
  assign _T_153 = {{30'd0}, _T_152}; // @[PEAlter.scala 20:26:@112.6]
  assign tmp_1 = _T_148 ? _T_153 : 194'h0; // @[PEAlter.scala 19:28:@110.4]
  assign _T_154 = io_b[1]; // @[PEAlter.scala 19:15:@118.4]
  assign _T_158 = _GEN_32 << 1'h1; // @[PEAlter.scala 20:34:@121.6]
  assign _GEN_34 = {{30'd0}, _T_158}; // @[PEAlter.scala 20:26:@122.6]
  assign _T_159 = tmp_1 ^ _GEN_34; // @[PEAlter.scala 20:26:@122.6]
  assign tmp_2 = _T_154 ? _T_159 : tmp_1; // @[PEAlter.scala 19:28:@120.4]
  assign _T_160 = io_b[2]; // @[PEAlter.scala 19:15:@128.4]
  assign _GEN_35 = {{3'd0}, io_a}; // @[PEAlter.scala 20:34:@131.6]
  assign _T_164 = _GEN_35 << 2'h2; // @[PEAlter.scala 20:34:@131.6]
  assign _GEN_36 = {{28'd0}, _T_164}; // @[PEAlter.scala 20:26:@132.6]
  assign _T_165 = tmp_2 ^ _GEN_36; // @[PEAlter.scala 20:26:@132.6]
  assign tmp_3 = _T_160 ? _T_165 : tmp_2; // @[PEAlter.scala 19:28:@130.4]
  assign _T_166 = io_b[3]; // @[PEAlter.scala 19:15:@138.4]
  assign _T_170 = _GEN_35 << 2'h3; // @[PEAlter.scala 20:34:@141.6]
  assign _GEN_38 = {{28'd0}, _T_170}; // @[PEAlter.scala 20:26:@142.6]
  assign _T_171 = tmp_3 ^ _GEN_38; // @[PEAlter.scala 20:26:@142.6]
  assign tmp_4 = _T_166 ? _T_171 : tmp_3; // @[PEAlter.scala 19:28:@140.4]
  assign _T_172 = io_b[4]; // @[PEAlter.scala 19:15:@148.4]
  assign _GEN_39 = {{7'd0}, io_a}; // @[PEAlter.scala 20:34:@151.6]
  assign _T_176 = _GEN_39 << 3'h4; // @[PEAlter.scala 20:34:@151.6]
  assign _GEN_40 = {{24'd0}, _T_176}; // @[PEAlter.scala 20:26:@152.6]
  assign _T_177 = tmp_4 ^ _GEN_40; // @[PEAlter.scala 20:26:@152.6]
  assign tmp_5 = _T_172 ? _T_177 : tmp_4; // @[PEAlter.scala 19:28:@150.4]
  assign _T_178 = io_b[5]; // @[PEAlter.scala 19:15:@158.4]
  assign _T_182 = _GEN_39 << 3'h5; // @[PEAlter.scala 20:34:@161.6]
  assign _GEN_42 = {{24'd0}, _T_182}; // @[PEAlter.scala 20:26:@162.6]
  assign _T_183 = tmp_5 ^ _GEN_42; // @[PEAlter.scala 20:26:@162.6]
  assign tmp_6 = _T_178 ? _T_183 : tmp_5; // @[PEAlter.scala 19:28:@160.4]
  assign _T_184 = io_b[6]; // @[PEAlter.scala 19:15:@168.4]
  assign _T_188 = _GEN_39 << 3'h6; // @[PEAlter.scala 20:34:@171.6]
  assign _GEN_44 = {{24'd0}, _T_188}; // @[PEAlter.scala 20:26:@172.6]
  assign _T_189 = tmp_6 ^ _GEN_44; // @[PEAlter.scala 20:26:@172.6]
  assign tmp_7 = _T_184 ? _T_189 : tmp_6; // @[PEAlter.scala 19:28:@170.4]
  assign _T_190 = io_b[7]; // @[PEAlter.scala 19:15:@178.4]
  assign _T_194 = _GEN_39 << 3'h7; // @[PEAlter.scala 20:34:@181.6]
  assign _GEN_46 = {{24'd0}, _T_194}; // @[PEAlter.scala 20:26:@182.6]
  assign _T_195 = tmp_7 ^ _GEN_46; // @[PEAlter.scala 20:26:@182.6]
  assign tmp_8 = _T_190 ? _T_195 : tmp_7; // @[PEAlter.scala 19:28:@180.4]
  assign _T_196 = io_b[8]; // @[PEAlter.scala 19:15:@188.4]
  assign _GEN_47 = {{15'd0}, io_a}; // @[PEAlter.scala 20:34:@191.6]
  assign _T_200 = _GEN_47 << 4'h8; // @[PEAlter.scala 20:34:@191.6]
  assign _GEN_48 = {{16'd0}, _T_200}; // @[PEAlter.scala 20:26:@192.6]
  assign _T_201 = tmp_8 ^ _GEN_48; // @[PEAlter.scala 20:26:@192.6]
  assign tmp_9 = _T_196 ? _T_201 : tmp_8; // @[PEAlter.scala 19:28:@190.4]
  assign _T_202 = io_b[9]; // @[PEAlter.scala 19:15:@198.4]
  assign _T_206 = _GEN_47 << 4'h9; // @[PEAlter.scala 20:34:@201.6]
  assign _GEN_50 = {{16'd0}, _T_206}; // @[PEAlter.scala 20:26:@202.6]
  assign _T_207 = tmp_9 ^ _GEN_50; // @[PEAlter.scala 20:26:@202.6]
  assign tmp_10 = _T_202 ? _T_207 : tmp_9; // @[PEAlter.scala 19:28:@200.4]
  assign _T_208 = io_b[10]; // @[PEAlter.scala 19:15:@208.4]
  assign _T_212 = _GEN_47 << 4'ha; // @[PEAlter.scala 20:34:@211.6]
  assign _GEN_52 = {{16'd0}, _T_212}; // @[PEAlter.scala 20:26:@212.6]
  assign _T_213 = tmp_10 ^ _GEN_52; // @[PEAlter.scala 20:26:@212.6]
  assign tmp_11 = _T_208 ? _T_213 : tmp_10; // @[PEAlter.scala 19:28:@210.4]
  assign _T_214 = io_b[11]; // @[PEAlter.scala 19:15:@218.4]
  assign _T_218 = _GEN_47 << 4'hb; // @[PEAlter.scala 20:34:@221.6]
  assign _GEN_54 = {{16'd0}, _T_218}; // @[PEAlter.scala 20:26:@222.6]
  assign _T_219 = tmp_11 ^ _GEN_54; // @[PEAlter.scala 20:26:@222.6]
  assign tmp_12 = _T_214 ? _T_219 : tmp_11; // @[PEAlter.scala 19:28:@220.4]
  assign _T_220 = io_b[12]; // @[PEAlter.scala 19:15:@228.4]
  assign _T_224 = _GEN_47 << 4'hc; // @[PEAlter.scala 20:34:@231.6]
  assign _GEN_56 = {{16'd0}, _T_224}; // @[PEAlter.scala 20:26:@232.6]
  assign _T_225 = tmp_12 ^ _GEN_56; // @[PEAlter.scala 20:26:@232.6]
  assign tmp_13 = _T_220 ? _T_225 : tmp_12; // @[PEAlter.scala 19:28:@230.4]
  assign _T_226 = io_b[13]; // @[PEAlter.scala 19:15:@238.4]
  assign _T_230 = _GEN_47 << 4'hd; // @[PEAlter.scala 20:34:@241.6]
  assign _GEN_58 = {{16'd0}, _T_230}; // @[PEAlter.scala 20:26:@242.6]
  assign _T_231 = tmp_13 ^ _GEN_58; // @[PEAlter.scala 20:26:@242.6]
  assign tmp_14 = _T_226 ? _T_231 : tmp_13; // @[PEAlter.scala 19:28:@240.4]
  assign _T_232 = io_b[14]; // @[PEAlter.scala 19:15:@248.4]
  assign _T_236 = _GEN_47 << 4'he; // @[PEAlter.scala 20:34:@251.6]
  assign _GEN_60 = {{16'd0}, _T_236}; // @[PEAlter.scala 20:26:@252.6]
  assign _T_237 = tmp_14 ^ _GEN_60; // @[PEAlter.scala 20:26:@252.6]
  assign tmp_15 = _T_232 ? _T_237 : tmp_14; // @[PEAlter.scala 19:28:@250.4]
  assign _T_238 = io_b[15]; // @[PEAlter.scala 19:15:@258.4]
  assign _T_242 = _GEN_47 << 4'hf; // @[PEAlter.scala 20:34:@261.6]
  assign _GEN_62 = {{16'd0}, _T_242}; // @[PEAlter.scala 20:26:@262.6]
  assign _T_243 = tmp_15 ^ _GEN_62; // @[PEAlter.scala 20:26:@262.6]
  assign tmp_16 = _T_238 ? _T_243 : tmp_15; // @[PEAlter.scala 19:28:@260.4]
  assign _T_244 = io_b[16]; // @[PEAlter.scala 19:15:@268.4]
  assign _GEN_63 = {{31'd0}, io_a}; // @[PEAlter.scala 20:34:@271.6]
  assign _T_248 = _GEN_63 << 5'h10; // @[PEAlter.scala 20:34:@271.6]
  assign _T_249 = tmp_16 ^ _T_248; // @[PEAlter.scala 20:26:@272.6]
  assign tmp_17 = _T_244 ? _T_249 : tmp_16; // @[PEAlter.scala 19:28:@270.4]
  assign _T_250 = io_b[17]; // @[PEAlter.scala 19:15:@278.4]
  assign _T_254 = _GEN_63 << 5'h11; // @[PEAlter.scala 20:34:@281.6]
  assign _T_255 = tmp_17 ^ _T_254; // @[PEAlter.scala 20:26:@282.6]
  assign tmp_18 = _T_250 ? _T_255 : tmp_17; // @[PEAlter.scala 19:28:@280.4]
  assign _T_256 = io_b[18]; // @[PEAlter.scala 19:15:@288.4]
  assign _T_260 = _GEN_63 << 5'h12; // @[PEAlter.scala 20:34:@291.6]
  assign _T_261 = tmp_18 ^ _T_260; // @[PEAlter.scala 20:26:@292.6]
  assign tmp_19 = _T_256 ? _T_261 : tmp_18; // @[PEAlter.scala 19:28:@290.4]
  assign _T_262 = io_b[19]; // @[PEAlter.scala 19:15:@298.4]
  assign _T_266 = _GEN_63 << 5'h13; // @[PEAlter.scala 20:34:@301.6]
  assign _T_267 = tmp_19 ^ _T_266; // @[PEAlter.scala 20:26:@302.6]
  assign tmp_20 = _T_262 ? _T_267 : tmp_19; // @[PEAlter.scala 19:28:@300.4]
  assign _T_268 = io_b[20]; // @[PEAlter.scala 19:15:@308.4]
  assign _T_272 = _GEN_63 << 5'h14; // @[PEAlter.scala 20:34:@311.6]
  assign _T_273 = tmp_20 ^ _T_272; // @[PEAlter.scala 20:26:@312.6]
  assign tmp_21 = _T_268 ? _T_273 : tmp_20; // @[PEAlter.scala 19:28:@310.4]
  assign _T_274 = io_b[21]; // @[PEAlter.scala 19:15:@318.4]
  assign _T_278 = _GEN_63 << 5'h15; // @[PEAlter.scala 20:34:@321.6]
  assign _T_279 = tmp_21 ^ _T_278; // @[PEAlter.scala 20:26:@322.6]
  assign tmp_22 = _T_274 ? _T_279 : tmp_21; // @[PEAlter.scala 19:28:@320.4]
  assign _T_280 = io_b[22]; // @[PEAlter.scala 19:15:@328.4]
  assign _T_284 = _GEN_63 << 5'h16; // @[PEAlter.scala 20:34:@331.6]
  assign _T_285 = tmp_22 ^ _T_284; // @[PEAlter.scala 20:26:@332.6]
  assign tmp_23 = _T_280 ? _T_285 : tmp_22; // @[PEAlter.scala 19:28:@330.4]
  assign _T_286 = io_b[23]; // @[PEAlter.scala 19:15:@338.4]
  assign _T_290 = _GEN_63 << 5'h17; // @[PEAlter.scala 20:34:@341.6]
  assign _T_291 = tmp_23 ^ _T_290; // @[PEAlter.scala 20:26:@342.6]
  assign tmp_24 = _T_286 ? _T_291 : tmp_23; // @[PEAlter.scala 19:28:@340.4]
  assign _T_292 = io_b[24]; // @[PEAlter.scala 19:15:@348.4]
  assign _T_296 = _GEN_63 << 5'h18; // @[PEAlter.scala 20:34:@351.6]
  assign _T_297 = tmp_24 ^ _T_296; // @[PEAlter.scala 20:26:@352.6]
  assign tmp_25 = _T_292 ? _T_297 : tmp_24; // @[PEAlter.scala 19:28:@350.4]
  assign _T_298 = io_b[25]; // @[PEAlter.scala 19:15:@358.4]
  assign _T_302 = _GEN_63 << 5'h19; // @[PEAlter.scala 20:34:@361.6]
  assign _T_303 = tmp_25 ^ _T_302; // @[PEAlter.scala 20:26:@362.6]
  assign tmp_26 = _T_298 ? _T_303 : tmp_25; // @[PEAlter.scala 19:28:@360.4]
  assign _T_304 = io_b[26]; // @[PEAlter.scala 19:15:@368.4]
  assign _T_308 = _GEN_63 << 5'h1a; // @[PEAlter.scala 20:34:@371.6]
  assign _T_309 = tmp_26 ^ _T_308; // @[PEAlter.scala 20:26:@372.6]
  assign tmp_27 = _T_304 ? _T_309 : tmp_26; // @[PEAlter.scala 19:28:@370.4]
  assign _T_310 = io_b[27]; // @[PEAlter.scala 19:15:@378.4]
  assign _T_314 = _GEN_63 << 5'h1b; // @[PEAlter.scala 20:34:@381.6]
  assign _T_315 = tmp_27 ^ _T_314; // @[PEAlter.scala 20:26:@382.6]
  assign tmp_28 = _T_310 ? _T_315 : tmp_27; // @[PEAlter.scala 19:28:@380.4]
  assign _T_316 = io_b[28]; // @[PEAlter.scala 19:15:@388.4]
  assign _T_320 = _GEN_63 << 5'h1c; // @[PEAlter.scala 20:34:@391.6]
  assign _T_321 = tmp_28 ^ _T_320; // @[PEAlter.scala 20:26:@392.6]
  assign tmp_29 = _T_316 ? _T_321 : tmp_28; // @[PEAlter.scala 19:28:@390.4]
  assign _T_322 = io_b[29]; // @[PEAlter.scala 19:15:@398.4]
  assign _T_326 = _GEN_63 << 5'h1d; // @[PEAlter.scala 20:34:@401.6]
  assign _T_327 = tmp_29 ^ _T_326; // @[PEAlter.scala 20:26:@402.6]
  assign tmp_30 = _T_322 ? _T_327 : tmp_29; // @[PEAlter.scala 19:28:@400.4]
  assign _T_328 = io_b[30]; // @[PEAlter.scala 19:15:@408.4]
  assign _T_332 = _GEN_63 << 5'h1e; // @[PEAlter.scala 20:34:@411.6]
  assign _T_333 = tmp_30 ^ _T_332; // @[PEAlter.scala 20:26:@412.6]
  assign tmp_31 = _T_328 ? _T_333 : tmp_30; // @[PEAlter.scala 19:28:@410.4]
  assign _T_334 = io_b[31]; // @[PEAlter.scala 19:15:@418.4]
  assign _T_338 = _GEN_63 << 5'h1f; // @[PEAlter.scala 20:34:@421.6]
  assign _T_339 = tmp_31 ^ _T_338; // @[PEAlter.scala 20:26:@422.6]
  assign io_pout = _T_334 ? _T_339 : tmp_31; // @[PEAlter.scala 25:11:@428.4]
endmodule
module PEAlter( // @[:@430.2]
  input          clock, // @[:@431.4]
  input          reset, // @[:@432.4]
  input  [162:0] io_a, // @[:@433.4]
  input  [162:0] io_p, // @[:@433.4]
  input  [31:0]  io_bi, // @[:@433.4]
  output [162:0] io_pout // @[:@433.4]
);
  wire [162:0] FMul_io_a; // @[PEAlter.scala 30:19:@436.4]
  wire [31:0] FMul_io_b; // @[PEAlter.scala 30:19:@436.4]
  wire [193:0] FMul_io_pout; // @[PEAlter.scala 30:19:@436.4]
  wire [225:0] _GEN_0; // @[PEAlter.scala 44:21:@435.4]
  wire [225:0] _T_14; // @[PEAlter.scala 44:21:@435.4]
  wire [225:0] _GEN_1; // @[PEAlter.scala 44:36:@441.4]
  wire [225:0] ptmp1; // @[PEAlter.scala 44:36:@441.4]
  wire [225:0] ptmp2; // @[PEAlter.scala 45:21:@442.4]
  wire [288:0] _GEN_2; // @[PEAlter.scala 46:22:@443.4]
  wire [288:0] _T_17; // @[PEAlter.scala 46:22:@443.4]
  wire [288:0] _T_19; // @[PEAlter.scala 46:40:@444.4]
  wire [288:0] _T_20; // @[PEAlter.scala 46:31:@445.4]
  wire [288:0] _T_22; // @[PEAlter.scala 46:58:@446.4]
  wire [288:0] _T_23; // @[PEAlter.scala 46:49:@447.4]
  wire [288:0] _T_25; // @[PEAlter.scala 46:76:@448.4]
  wire [288:0] ptmp3; // @[PEAlter.scala 46:67:@449.4]
  wire [288:0] pGuess; // @[PEAlter.scala 47:22:@450.4]
  wire [543:0] _GEN_6; // @[PEAlter.scala 48:32:@451.4]
  wire [543:0] _T_28; // @[PEAlter.scala 48:32:@451.4]
  wire [295:0] _GEN_7; // @[PEAlter.scala 48:52:@452.4]
  wire [295:0] _T_30; // @[PEAlter.scala 48:52:@452.4]
  wire [543:0] _GEN_8; // @[PEAlter.scala 48:42:@453.4]
  wire [543:0] _T_31; // @[PEAlter.scala 48:42:@453.4]
  wire [295:0] _T_33; // @[PEAlter.scala 48:70:@454.4]
  wire [543:0] _GEN_10; // @[PEAlter.scala 48:60:@455.4]
  wire [543:0] _T_34; // @[PEAlter.scala 48:60:@455.4]
  wire [291:0] _GEN_11; // @[PEAlter.scala 48:88:@456.4]
  wire [291:0] _T_36; // @[PEAlter.scala 48:88:@456.4]
  wire [543:0] _GEN_12; // @[PEAlter.scala 48:78:@457.4]
  wire [543:0] _T_37; // @[PEAlter.scala 48:78:@457.4]
  wire [543:0] _T_38; // @[PEAlter.scala 48:96:@458.4]
  wire [543:0] _GEN_14; // @[PEAlter.scala 48:21:@459.4]
  wire [543:0] ptmp4; // @[PEAlter.scala 48:21:@459.4]
  wire  _T_39; // @[PEAlter.scala 49:23:@460.4]
  wire [162:0] _T_42; // @[PEAlter.scala 49:43:@462.4]
  wire [162:0] _T_44; // @[PEAlter.scala 49:51:@463.4]
  wire [543:0] _T_45; // @[PEAlter.scala 49:17:@464.4]
  FMul FMul ( // @[PEAlter.scala 30:19:@436.4]
    .io_a(FMul_io_a),
    .io_b(FMul_io_b),
    .io_pout(FMul_io_pout)
  );
  assign _GEN_0 = {{63'd0}, io_p}; // @[PEAlter.scala 44:21:@435.4]
  assign _T_14 = _GEN_0 << 6'h20; // @[PEAlter.scala 44:21:@435.4]
  assign _GEN_1 = {{32'd0}, FMul_io_pout}; // @[PEAlter.scala 44:36:@441.4]
  assign ptmp1 = _T_14 ^ _GEN_1; // @[PEAlter.scala 44:36:@441.4]
  assign ptmp2 = ptmp1 >> 8'ha1; // @[PEAlter.scala 45:21:@442.4]
  assign _GEN_2 = {{63'd0}, ptmp2}; // @[PEAlter.scala 46:22:@443.4]
  assign _T_17 = _GEN_2 << 6'h23; // @[PEAlter.scala 46:22:@443.4]
  assign _T_19 = _GEN_2 << 6'h26; // @[PEAlter.scala 46:40:@444.4]
  assign _T_20 = _T_17 ^ _T_19; // @[PEAlter.scala 46:31:@445.4]
  assign _T_22 = _GEN_2 << 6'h29; // @[PEAlter.scala 46:58:@446.4]
  assign _T_23 = _T_20 ^ _T_22; // @[PEAlter.scala 46:49:@447.4]
  assign _T_25 = _GEN_2 << 6'h2a; // @[PEAlter.scala 46:76:@448.4]
  assign ptmp3 = _T_23 ^ _T_25; // @[PEAlter.scala 46:67:@449.4]
  assign pGuess = ptmp3 >> 6'h25; // @[PEAlter.scala 47:22:@450.4]
  assign _GEN_6 = {{255'd0}, pGuess}; // @[PEAlter.scala 48:32:@451.4]
  assign _T_28 = _GEN_6 << 8'ha3; // @[PEAlter.scala 48:32:@451.4]
  assign _GEN_7 = {{7'd0}, pGuess}; // @[PEAlter.scala 48:52:@452.4]
  assign _T_30 = _GEN_7 << 3'h7; // @[PEAlter.scala 48:52:@452.4]
  assign _GEN_8 = {{248'd0}, _T_30}; // @[PEAlter.scala 48:42:@453.4]
  assign _T_31 = _T_28 ^ _GEN_8; // @[PEAlter.scala 48:42:@453.4]
  assign _T_33 = _GEN_7 << 3'h6; // @[PEAlter.scala 48:70:@454.4]
  assign _GEN_10 = {{248'd0}, _T_33}; // @[PEAlter.scala 48:60:@455.4]
  assign _T_34 = _T_31 ^ _GEN_10; // @[PEAlter.scala 48:60:@455.4]
  assign _GEN_11 = {{3'd0}, pGuess}; // @[PEAlter.scala 48:88:@456.4]
  assign _T_36 = _GEN_11 << 2'h3; // @[PEAlter.scala 48:88:@456.4]
  assign _GEN_12 = {{252'd0}, _T_36}; // @[PEAlter.scala 48:78:@457.4]
  assign _T_37 = _T_34 ^ _GEN_12; // @[PEAlter.scala 48:78:@457.4]
  assign _T_38 = _T_37 ^ _GEN_6; // @[PEAlter.scala 48:96:@458.4]
  assign _GEN_14 = {{318'd0}, ptmp1}; // @[PEAlter.scala 48:21:@459.4]
  assign ptmp4 = _GEN_14 ^ _T_38; // @[PEAlter.scala 48:21:@459.4]
  assign _T_39 = ptmp4[163]; // @[PEAlter.scala 49:23:@460.4]
  assign _T_42 = ptmp4[162:0]; // @[PEAlter.scala 49:43:@462.4]
  assign _T_44 = _T_42 ^ 163'hc9; // @[PEAlter.scala 49:51:@463.4]
  assign _T_45 = _T_39 ? {{381'd0}, _T_44} : ptmp4; // @[PEAlter.scala 49:17:@464.4]
  assign io_pout = _T_45[162:0]; // @[PEAlter.scala 49:11:@465.4]
  assign FMul_io_a = io_a; // @[PEAlter.scala 31:12:@439.4]
  assign FMul_io_b = io_bi; // @[PEAlter.scala 32:12:@440.4]
endmodule
